��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����0� ����遼�6������"���#�{A���'j�Qj} �}xT	g��F����a��f��洜K%g==�Z���L1������bG����XB�k6T��w+F��3r1#�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf^��$�i�g�Wɐ�)
�Ql�Y�+6�iѰ�^���d�u�.�Ye�ZG�$*�f�pM��Y���f<���YB�H6]��^�8�G{��:RjeQ��2
�ƣː��5JLO%/.�)����\�
,��YIw_�aJ�/��]b<Q�	������*;Rdn�����nG�"M����u��~8�
�����a��E��{_ɸlw������e0�P���EY�2�΄��Y�n�?��6�$-D�T�%�[��\t,.��c��Ⱦd��ֶ�5�6}Fh�H�J�A5u��yOj+>���g��k���LG�wrث���)�Zm��toN|ٹG�Uk���4�X��;̰G*k2�bI�p�-}-z�Ń���KB�_2�~��j��7+3��PǇz�D�ˊܣ/D0P��4��i^��JȾ(L���5�iF��ӭ��c@ܳx���	8 ;�5��_%���R��gP܏�Z�lW2��p��/�)�tpR-�?d�(?�(`q��r�Aͼ=��邐�|L�}nx��osz��>��<��*�+��tU�;�{8�r�{�d�eQ[f���4�V�	]��"�h1Ӣ'�g$��91���+�2�=6A�(T�sl�l!�}�Q���|r�����Z�;�5���O�D/�im��+���ji.qԞ���}�"��q�8PX�%]�&�e���6���%�h�\���>dL&ї4U$h:�0 $�l%�`��m�� ;�6���'.�'֛c��n�Ǟ-L�R��ŏ����2U�e����� >_$�c�>�C��k�5<��Ş�h�ݺUw�p�=�k�\��|ot�m��}r���]�:ܑ��J|n�4�i��1�|�Vmc<b8�u�3eu�U�3,�Q�PM�K�w<�2����0���vN����'VlC<�ap,9י�ч�D
J�I�2J�M��dK��:��rjS����^&�h�09�(Z�n�!�%nz 1�kkH��\��]���X��+Yh;p�:#��imY[ý�嫃�ƴR��e�D�_W]b�L�&T/�*Κ����߿;1���# ��z'�ؤ�8{*�&&�靽�'N��z�K�RK�y����ϭ� �@����g3�7"��r��*�j~N�f�[�Qe_��F*3.8��᧾����ٮw8�1ΨκB ��X����m��f�'�lҼ�1[N�s����A������R@+{��&�ѐT� Y��x$��/�0�j�7{�Ճ�wex�"���)��'gfv�H�b�@��P'�����
�4ki+2|/Qm�	�v���xK����E[է��P �ֽ��t"�%Vb��,2�Q���t����$��@y���qH�F@�ӚP�߫m��đ��b�g%�$�oD�B��
C�S�8�U@� K�b���Qp�<x����}�����y���3I�!��8>2e?*K�x����r�>�����S���^��i��c�5 ��q���/O2NeB�X�ƃ�?&
�7��Ϗ��|o|�j��_ըY$��Q�ǔk�Ɣc	b��6���_��i����5:b���v�X��*DJm�yh7��i�D�\����2�,��R ��+2�h?��>�r�:�Z:t�(����F�e���"�n�F��ˊ������V\8�ϒ�lC�*�pݿ��Ӵ؇���N��N�H����3���2��$ә�⡲�!.V�����O�}� 'RQ�>Y��Ov�Tj8��nĲJ��6P�.?I5���=�ů��������-��j���ü:C}�8+��/uun���tcՅZ��x%�˾���}̐`uw#���*Պ,/Һo�r����dq�6|/
73.�m�0���zboP+��Bn��O�u����h��e4��r����X�K�7�r���R��W ����M֞sը�9�<X�G7*�g�;����ЙQ�s����(��N�ݺ~�����?K�6{��1��*��~3��=L�c��N�G��"ϰ��*(�݊4eH)v��l�?x�h��`t�g��l�ɟ́�␾j%�:p�,��r3ť�x�w�R#��վ�J�|�9���� U�:ڦ�!���A��* ���
d#0F���Ⅻ���?[
D����s�@�<!>��+�B=��_��ԧy�A�=Va�K�ֶ�ҥRm{�ȵc��D��W�}0��°a����e�5_�70n�����Xϵ����W���<�р��h�,�G�dC�y\,a/m�f��QI����#r\�YBtK �n��f�P��I�[|2^q�]5��SQc��&��:�$�<k���{-�_�N�u�� �R�G��Wm����l�	�䒴=��8 E��Vn�)�D�ܯt9�{�8�;z�!T�Z�j�z������� r�����Hvh ��;i�t�֖&�g;h�E�K�'b��k���8�'�?8щ�����Ut5�S��M�cx�`�#8.���q�[���)��}�sb��{­��4�c��ݏ��t���.�����헆�ӎ��:�X�֕tJ10g`9V��84�D��wj��>��Ĕsy�S49�!���ȩ?�-�(_:L!07v���Ǐ�G�m6�^�2�������!l�Z��Tlǐ���F\�8�6���9��휆̍�8?��%X���C����M�_f����枭�]8���0��g�Riy��/~@��g�nעxD�����^����V����˾����p����W�6!��:,n+!� ��di9U0Q�ht�9���xq�c~�����	Ǿ�QI��M�Ѹ˰�`� �m��˨Km��3���I���&fa�-�1��w�ٗk& `F�n;~���\C>�S���'p����J�6��"��/�-4�<�}-d�#���)�Z�I}�ḱ���K��׻cg�"N���CM҄В�x� ۵��\,�H��'M�Ҳ+[M_&���(S:�`�L�X�<5��!�>�q��0IvPE*od�=1f�&�WA���5�r�%nX�pҞ|�XEV}��A��Q�i7���C����V�	���0ɓ���Kg�'��m�E�=S%���s��fLch������P���qꆽhA���W���~=a�s������I�术>������Ϭ3���dt<���L;��� ݨ��,�d��P�E�}��\ȶ�C_yzV��QM&�����5���N���m)=n�7"E����q��e�5��`�	���%�P��/|���Iб�����;I��{�BΤ4����+/�a���š��=6��o(������`IW���S�\�Zf�Jm��������BE�B��A��N@��^ݼ��}��@���Ud���))��&��d̷u�%���}2��W�qP��ZaՓ�5�����j�N ���;��;Ҹ'+)O�re��������ǖ&��VZJ[�Z�A!cn*��4 x���CBX&@����/8A�׽ą 3��*�o�n{�,�w�zw���ٵ\0Nݱ����
F���!�N��;�e��M~	Q���*�>��h���=N<�!�zʣ���B�4x�<��!���x�&�|��m�ʃ�*�t��->�i�����7F' �?.�_���R���0� ��}�X�u�����^��Nh�W���]1cr�D�� %��$���o�i*�l
��-�S�ƪ�D9�U[UVWt� ���`���߁��g��,p	���������>A*+�w<[�7����$ ��:��
�<��$N}")X�SMh��y���oTl2�b�Wf��0�/P��+¬:˦��	�F��$���1���~��_��2����"u�K7��S�7�ʎ�6(;#v�s*Rk:e�9ͪ��Ra��Ve|i£�.��QJl�N����bz�&ӫF���"�?OY�Y�kX�E��?3�=-X�rF�ҵ�*w�vw��Ђ5�hQYvD��q�����h��s��E��:��n79�$�R�r(n��.�����@�"�������5Bv!I��0���x�^�������n�h�f��@��s؊<Q.FŁ����^��y������*����'ۏw�G����d�n9�u�0���Q��у����|2:�;�Np�==
���|S���1��w�g�����4��I�|�H:Uf�����Z �y���M�ڝi���bM���~���7��13<��)���"qT�JX`��Z 	�osR���k��jF���7D�ヰ��S%z� [��n�(bzڐ�f�h�*AF.&��=;a�>գ╾�r$��)U~�Ч�,���4U�E}��ǘAbN�6o�����-wΧ��=ƙ3R��	�|�i�e�T���p`�Oj��b��|�εHUO�S����W��(^�����H	��B�b���Pg!6���r>4\���DWdk?Ҭ��6��{�����# �;'i���QR�4�� ��f�j��f_�~��%æ����9BkT;xŲ �e��SV��3�V���i4h^��c�!Q�R�wwd�\�o�2j���q�g�b���v��8��;�u��y�ӗJp�ܒN�R8�&�?�������*�2�D�Yvpm�@�v���F�Sl���}�y���a����Yg4]�H[K�4o�ݔ�&�_�?���V���.����GX��ܜ��)>�%�#]m2�%t{�30���J`a�$0��X��߬_שW��0�.Pm.��%?Ԯ�{�/.*��F�N�=\���+�xX��� hm�D���&��.�kW�UJ����֫����"B�����0�JV`�t��/��c_����t�W��������b�:k���Gt��y���r�?���>I���X�"�?X�Pg���E�q�r霬���'ݽLU���kj���ɄjI���fhk,H/�h���Ul����@���5�)�19G�	��C��->ġ i?o_`w�=�Q�i�-I��S��ۭ�X��vJ#:��/�������p�X�-������ե��L�eC�D������,Be��SPP!X�ԁ"�Z8�8������ D�4�0�O�t���"�ZE�~�+�h��7G�"�5��DPR�cD*�F^��_k�%)�h���o����!�3(��>5&�e ���p�8����.���Nh8����[l:��%��ld�Ͽ�V�|���X�=�J��8C��DH!���5V>s륇��w�=�ԥ���0�h���i�XK1Ba�)��Q�f`Ŧ���r0V'�V�Mi��F��tD���hg_c����C��[7@���B4��{!XJEJ�j۹K�����N�VgL]��_�<���������}�h\��z��I����R*i���V������K��g�3}�����;�d����A�stA��w��l��*�g��v*f�ɯ��Y3��'~��ɺ���l͖e�;U���dȂ	z;"u 5���m�#�M&���2 y{�1'\��Cd\32�DA>JK��}
D���/XFG�+˫�g�Ҵ�T������*/~o�V'��ȫ�5�Ng���Y��(nŮ:W�.L�}����a��r��p;ٿ�K�*x��2�C�����B�`\�.C�h���|�"1:�_ۻO~��id!Ff�l��8�П�Ky7x#I �@`OW��6Nm%�����g�*�!0bOP��
�<�c��qBGtb���t�cK��S����P�����&u�I�S��(�1����
��::�g#G��l�����`%L(!�4�����RwIJ�|Ju8��l e��L&ޚ�wMM%T��m�m��x���H��K<o��	�G�͛�ă%~�h'�dnl�1aƯ�pB�X�a���>�eB������#Hg�:���m�ٔ��3�'zI�`��Oׁ���e��z�}�W�����>�� y��/��Z�c*���]��V*�4kU�)�\�;��%���*�ga��:�������s�ȭ)07���E���9��O~��i�e#�OV:��CK��1��C�5��dr������� �Mk�Ue���)̀M�N
3�#.���9� ��$Oyk�7$gU��
��)�5���iL:��l�i�q%9L�չ���d`�)�x�]�y�/�1����'�����ل��+�41䑹��X��j�Tb��P"�����{/6,���s�M�.C��USV�D8�K3���v �H1zP�MK��`�w
��m1�О6�n��#�a+��V
GaS��a��h��ɉq����׈]l>��ȴ����M�9��p��j%�o:�s���(�XZb�6��\��Yb5u��'�إT�j�)&I���ϑ�b�A@�p��@b�ӛ�`�@뗖���^q������}4�d�!Zj#�WM��ZY.	�Y���pH]��j��Aq����\q8m`�+Dr�y���3�h��~�v�_�$��H�G����|}��N�b��/N�ʌ�b��>y/Mg)��{�	�)���J���'�ٱ�G'��*1�U�I��O!p�r����<�.K��#�>��흆�D�}B>���ՈS"y-#}���xu>qAo��V�u�,�7K�IF�˘�S�9N��vy����9a�^���S�W�����$2OZ�!dT�dg�q�BТ;�? ���p��ة��s��t:���0NV^6u	J�2���B8����j���*F��c��.���z�&�� Ry���ȠH)�l�E{�K�=,B������3�Q_t����<��o�'��� n�8���hyV^Q���jэ�q_�;J�$�|��gΗg(�o����Z�VmN���'/J�2�[
%Lҿ��n|�(�:���7IR8�$[)��*��~�� IZX-���X�3���p�x�\Q����f�Wj�M�X�*v}
��<S-�ϭp]���-8V�%�0s�ZOX[w/�G�((�I���X�^፵R��z�^�ITM��Oo��0O�uu9E�r�J�&�~�T���D��jq��}jrS�6����>A��Q7���I���m�VTPp�<�p�c�qx�j�,�[�������ӛ�(g��f��fN�KR\m��&�5�LKv��xi�0�!�����dyD�����w�ѭ=���
T�?�rt���Œ��
�ֵy�2�&K�O�g`q����rh|_0�W`�>�̽��$��
`�$C/NOr���Th��rӊ�$Q#(���,��E����ts?�xyh��^y
	ғ*(̋b��l*e�lf�FqȔT慒�8��5쵵�B
���tqo�Tk��lᒱ(��:�+�"��{_�F�Sf|�9ي��rŻS��0>Ja�3����UU[�|_#%���m���C�H�u���nXV�1%�5�"!u�u���F��}�@j�����۶��IO�GQ�rc�5%6~aq�� �&�H>nJ�0���>px�H
�����_ߴ 6���h���w��A� ]�.�{�/�S�!�gt���C�C,h7[� �k��Q�<�������n��"��km��$�(]�t~��ޙ���H$E�p
��s���<ZN^
��&��ya�$��!F�19{�t�}��iO�13�έ&�^��.����B���i�r�T4���D@�m)u���l �]�Z�^_����5k?�y,T=<s/��!���3�#v�0c�/�
|�ݞ%�+'j���p�kk���.��� ��� pb�:��9*0\��/��{� ���^�7~�q�)�qPe0Ѝa��3$o~�����{�5��>ZQ//723��6'�bo���U�����:BY`�&��~��͢�<n��"��R��|�������˄+y\�������+���vȄ#x�>2�:���Kf�������ia<�����ݫ ��م��D�$��G0_�r:r�aDR�-��>�1+�+��o�(׿�;�/�B�ԫ��LH���G���X'���7A��ˊ�PX2�?��X����b�� eH��=�#�8W�k���S'a��A�PDT9�c�C���+Ǿ�,
��eI>pn� EK���3���[��q#�����@��bU��6�1ջ'�A'ME&׿�s~�L�`.���.� h�;�J�ߌ�����/i�Prv��Ʀ.+1����<B�E�\�L���'q�ڏ�Ʋ��X�2�f���3/���c� ����B��d����t��<rއ��#r�����.���AY��J���b��yN7�.��_v{��u����I.�g�� :��xj�B��#��\���'�R �y�V񶲒l.���&�j�^��M�io��_�|�[[}�;�#������)�y��_Jj�s�ο�,�b#��Q!�fx�8���E,�G��شӞ	�Cr�*"s"!8qƛ���� ��z�;�����n�ۼ0�wŪt@���D����	�R�	)S�s�Q)��Y�,Z�Y�Дc��E���نYs� ح�㽻�P�[�<�@��+723Ʃ�S���H{�ƺe����� �)��Y�i{�p�c	Պ��J�H���!����.j̅�J���.7#��x�g+��7��ޒOcU����N��u|�4�@�2��*�J˭ITޔ��VX�[a�U57�7�O#$���q�����O�}�@U�X��z	�������(�LAY�37apN9ӌ��2�2�[�ʱ;<]�s�y���5���ϑ��/v
��j��xE>N�LL��A�\5�_q� �;�f��+��}Bp�+b"k��D��3���W.���,�UB�ϓ�j$ڐ��+�\���n�O��D�V��-i�T(�=�4��hі�	�_��i��cw44�v�a�;D'�^�� N��j����|Jx�^
t&̝Le�mɠ�&��E��cw��[��7���s��ut�s;&��,g��ľQJ������g�	��?k�b���|԰4!�"�� �qE���:�p���Ԅ_1<�E�e��9]��s2$�I�/�L�Z4~��ƣ���
��ͻFb�t�M	C��C�˰v3���M3�͝q_��V�L���y���!��0����b�<��E�zp@�~�wʻ��'!ǒ�B,y[�bX$��/�����=�0�W|��*�l�LJL��^�Yq�h:P��D� $���ww~J{���Y���o0��1"�&�y�T����%�3��R�c�b�t���Y	�S0�F��5
�T��/5�@��i '��$v�������{A&���l$����7slR��9�Ԯ�MlD}�+C��GM���~f���yI����yc���r;�B�´�PFeBǎ@��������42���"4�{EQ��is���!xx��G� ^_��c���"I�t��+dD��z��.�OC/(p�Mu���]�C�	Ԟܸ��f�=#�3�J^�>��z�'��h�SFr��Ɋ�;��P��g;tXj���ޢ��pֳo��S2]�'�)���%�E�ҐVu�{���'�f��B�{�jG譝i7ݠ��.��]��dd$�����6!y?�
X�1Ӽl���T�G:2r|�#s!p�y�(�Kg��f$(4޻��o��?�̓ܵ��>{��l��-罱"�0�2�v��u�Հ��ɳOu��%���*Ӟe���S�J������%s�����`�3�+Rkv�X1�#;Qd^���)�%���q���5�V8��������s�a��@��s�!R}������c������ڋ�D�yﱎu�{V?��7��4�`T-��)���_gw��V*����8�E�$ǫl��tI��]a�J�ؙP�V�x����[��a{�'�>z4���L���ڗQY>���J��;.ķ���%K�8 �k�<��*o9T�R���mf��	^͖�k�Z2��$��B�	��z���7�ڞLW�ߡbǇ^�S���A�I9Fs�2���
���x�ȁ�'�K.�|���"]j-�=�\�b�����>N��"Ee�őo��R�0��@��C�n��iȢ�Q��!�Z�!��=�D��'>�JN'�����q��=�=����~�VB�t2�D��qr
��׵���c������K�����
�"�R�2���˺7'� 4W��7�ÿ��<��E{_�N'��bW�cX+�b�P~��[鼧��z��S�K�3Y7����;u�7���T�v$�mf��@��&˵�"�#���q���8�x$NuǬ0*��#O��m��Byen䮫a��m��#��?3��C!���¬C�A�ޘ�O�q�����I͟�h�3�� �a�c��|�ŋ�6��e(���oYd$X��炳��T/����HwIaJ�$;4�!���l��>vݐ�'��A%�Y�4��_���y�tN��\ܒz������ �,硳h.UoI�H�_��9�u(��Ѯ;�^�Vz�1o 2��7�8�#�,{����q`d��|�H�Xu�qU3&"� 0Mq��)I�(�#� �GS���%�������S�]��F��aY�.b9Q�G�w����`aX�Lȱ�(�C(�9r賲F���{���.�u���u�<�������g�?2��Em��!� 1��_~�_���~��I���Փ��s�I`���B���:�{�������T� ����B̳��i°�)�]o� ���PL���؄�Ak<Ӏ4O
c�ħ�`�V����
��_P��J�����f�{���;N��{ ���� bt�߀qUW%٦+�ym���=��ׇc*#���[ٷ�[�x�:;�M�8�H'ެ�Mta�,��&���Sc�w�a�q�0��˂�3�-mTomX����SUͩp|�z
��s����>����Ĭ�HA�o�����Ѫ��{�ʅ��;z����+?S�v�¤)�3�.(%FSF%Fva��n��9}���P���~��+^>pFY�L�#����?����$�>4$�5)��ve��/p�SN�}(��W&H7��Y�h?��~��`I���a�!(�3�9�8�c��'r��TS]�Ի]�Y'�ϛJ$���]�nXU�<����zn,�M�u��h˸"/�vh��p�U���>6���q�;L�e+J�Q�{�ҕ�vߦ���U�5>瘈�-�YM�o �yޤ�ԴH=���U�4	՗�}U,�;��[��=	kFa���^l*���:$��2�n5��~�Q��B9=pd��Ғ���z�[j'�W�\�2N�[���#��A�&b��B)-�"T�Pa2Q��g�Y���5��X���%�$-Px*������o\�����{B;!�����~a��GP��7��{I/��\C��)��#ف)��� ֚��N��B�*�07ѣ�N��C�u��tv��c���z�CCxYϻ�
��Y�w�}o��ݑ�B���_<��mn�p��/��r\��r��PLƆ��g$u�`&��ʈRM�kW&!����E�Z�?�Tʜ��|pLw�~f����_|B���,j�h�>( ޟ��+{��ԁ&vUY8Gl���qY&�5��o�Ҥ��g���i��b�k�n�d�
i�e�J�����&	��1��w�������*�C�Py9� �Ɩ�7��ݻw�>WJ����A�����]������[�#a�2��ؐ��}XsזsN��.�A� ��]8�4�m��l�ǟ���J�r��$�Hv|M	Nv&�J���~�#����	��}�l���?\�.RaG�%f��J����+����hj؎Ʋٚ�4*fo�rΞ��:r]]�����J7Ζ#N�ho�J=�.FgZo�N>r�GN=W��y�����#��D<*�OQ�C�@{F��i�(N�.X��	\M�+9�"��lj~��E�w�C���.Q����pڝ�m���t9	{����=\�n{=_��8����_���Ё�d�(��.D���G�`����kӴ��h�J	�=������TK��G��M����7��ݰYH�g;U�r�r�ֿͲ�@���c���[�H��S���]�S^�"�v+�y�j?���^N��Ca@SM�����[w���J2�8���jbac����h����ݦї(z�eUw�1}IAe��c0@��/�1�*����d�1�g�T���4�!��r@P��)n�@H�]��IYx��t����k�%��#uV-���iN����-���a�g���zĊ�fc9ì;e�MC���|�C�d���AY����ף_����D�
���6ώ��~��C���W9�-\p�W�V��9P1��\��xd�G7
����"�V�y���	�� މ������O�D�?O��%3��)�֢���(#7] W��`�V�;P��4W=�\B�Zr%��B�ڳt:�����x����Q���Ά�`�H��h��l�Ԡ
����:6�RO���4��C-�/)JU>ez��S��md���.ǳ�F@��^o*�6܈�Z�YÙ*G�Ȧ�"|�� �r*KA z���L�T�9�Aw��+�)��ze��M�h��\5s�/���j#!��/��"Bc�ΐ����_�)�
@���4�R�vYMB�c�u��L������V6��|�'�?9{7��P���E�=)4�7��w��w��R�:紼��pe��|� "�!]�Mg��P]�ǡ���/��,�[۰��0��m�V�Kʄ�g�cX
��N�M��	���=�`a�ٲ�H�0��t�W�����'ń��jY�-�E�o�qc=iT���l�D��,���6w�d�`���䫋����H>�կTM�S$p��������1#9pώD:�e�}
ڨ�T������n��|xf�sS��Gf������>�3�_e��\}�Tim����Z��fN���k�2�V��S�z��)�g2���58˞U����!�?ŏ7�ۣ��^%�� N��e�k��������l5��mtq��"V�ġJ�.F�	�z-w�	Bt�t���w���^���P����q�)�96�'DM�C�����r���m_|h���*�꽕�(G&�Uo��a-,J �V2���'{䓦��N_U��ݦ���Qm�0⬲����f��М�@�i�g���2��q:	�W�I<RkB�8ٔʚ���-��C�"eW� W?#���%e�G��RRA�]���x0+����+�{�\�Y�y�Ѭ^֘�O��PW���1�{��q}X#�%�K� J�ޤަ8�W�/�j���䁒�E��� ��|&�^&���g�4=L�O[$=׆F�f�J�c�UN��ӱ��0o��}�W�03�Z��w���� ���i���)�|�.N�H�}٨44Bq��<�B �o�W�����`��e����a�j�[�.��ف���5_�'p�Ⓠ$S
؆n+���ć�E|���>��l��PehP/7��}�M��a&�L���_�}��t}4�_�uc�>��:��z���,�}=n������B\\�M����1��wKQ�iG&5����𶡶�~�k�} �4ӧ���N%��~���CM��9��Q�ygE�
��J·�U�l�QA'��<�D�6�w=9�Γ��ݤ����1z@�{A�D���n6�����8!�=ݼ��n|
ںf�����'G��ߖM��$��2S/Oz�0��*�R�G>�qLd��.+�������w���Q5��F�f��^!s��E$�ѣ��7���9���!�b`�76(u��|��Y�oġ$`��r��XJ1`��?��%y����.���?�ay~�� �ݙ_���_L�LX���^ŠϷ���� ]^N�@>�=>�١�t�F|Y>>���fa2�ؕ���L^����B�g��B��{�<�o�d.���^a�[��q$�D�R��?Si�B����wL]�5�J�Y�N��y�z��rr������tN��8�BX����bO	Q�sF�Ђ)Z��U�x�_�ZiF�w�t� �&fc$d�����C�CnQ#-5�x����
���'A{J����2ۄ�S�'�dX�Wo��E�[OU[J��#@"���	��1��Q�����@�5��3g�Z&�z��Y!=u�ݬ����6�<�|u��j�eJ�Հ3l�)#�Y�4gΰ��J�+oA�:�,d�����d�:�,`���A��F�QbID�ڌ�xf�����6���ñ��U?P�.��y�"���7w���ǫU�(>VM��L�PfG��Ɂ��=����wr�b���h9@��r�qͿ��FA"�2=Hiq�쾯���I��H��v��unp�cb'B��>�Y�jTu���qg�j&S#*%��6�x����<%?��ZyM�/34D��2a��[_~_����f�[��C`b����U�oƆ�Y˥3"z����X�/����d�h3�ڴ<�p V�_�꣑v����y�oORgߩ���'h�?�W#/�<��w���M�C�5)�ZVi��}�,��[��LRȅ�J5lr�v���Bʍ�i�*ۘ���/�o�kM��z�+�``s҈�&V�O���]owja^¥Ȅ�(=��
�2}����p�_{o82�e�qS��o,,���t'_������������:�� �N�\��v��p�P!g3pj܉>��RqO��:ȑ
u��]��q\�l����d�����`�'}���R0 -�d�~r?'B����s��$V���{�k�/q��*n�W��M�`��N�Hj��IRˍV����ϖ 6�b�SdRʈh�O��XR �I��!�qar%uI/��<�;=�Ķ1�m^�t.s�ϲ?��<�ܻ);+w�4��l��6v��	�W�����{����B"�9���\Y����Y�~z�b�U��h��I��`i�T�;[`Џk�[O����ٟ�pg�ra%���G�tb<���3?rh��2b�K�����y���m0?�OU���+nG�#��"��*
9�A�u�Q�1;��K)'�N��OA�Q�,I�5IW��4����=_D��e٤�N6�}tܱ�w���nT��K5�?O+ߋyj��OU)��d���#l�:���1\�ʫ8z���4>����G$iB�)�|T�w�ݰ�6�EX��7�	� �~��8𯑱�E��I��Kg4z�������(k�"�"�[Y~b-#G�|?�ɶo��.��WM�Æ�0kM�rѣ-���Y&N�:/�Qu�d�M�DP�ĝ��g,4��Kd����ǝxhE��쳞�A^��:z}��J�ҳ�`�J�b;��7f�a9zUv;D8KW, zÂ��f=�--s�Dz���R��
>�M4�q�T�9��;��ZE��N%��q{_6�(�n�YѨVF�¢Tօ���X��|�x�o+x0�v��D�>I�!�ai��&= ��ʫ�����/ڹm����E�<\�Un��`@V�� ��_�uI�p��#zJ�(����Vc�1�B�H��җW�4=������@)�n����E�4�{K��۸N���$����*'��Ñ���jxh��A��~���S[��׽#ӟ��ʘ��KEҰ���|�zk[��ޫ嶯���%�j6Zٮ����_� ��u/� 3:�"��L�<�`D���t�G�S�����w�G`��<3W��f�g}��$&��������.�1�8º�00n�"(xֺ�)M7^ћ��7/zfϏ�PL��7j��꧲�n�~��z���?Pk�FdK)�J�c�QF���v�9��O�-)1��D<w�rTUP)�F37�td�?���x�*@<��r��\�:����r�1^�� zh�(R��6rO�DUІ$�{����"��7O����S�'��M��)S�y����`��lP{6��j�;�����<y����_W���#���P��^r�����qEk�pr-Dì2y>�\Aѐ���ZL�.���|~��yJ3+��w$����=�^�}Q~�i�c��BJw�����5��q�e{�����Xu�6L�v`u�7�n+�6�4-�H������c�Q˗�ԅ����x�8;��Ɨt����u L�|g4�C�=g؜�?	4�Pে���~c�D��:�0	J
��l� �s�zU�&�H���fh�K\�X�~�ܖ̀?�l�󷺲;5y�>���"�r�a.�Rݣ1�_א�-�^1f���-��+�wXiH���S�/��Y�Z�ܸ.�!h�V��*[[J�;G"��@�3"��~%oQt)ni�$��)g����pj��I�iA?;4\Jt!��������R�R��~|����r(�G�EV����v��G�o�L�y�'u�x�A��qቬ���L��h��ZW��0�4�ܑ\�~$�FJ��5]�I2E��<	̖�Q�ā���m�ȅ\�Z"a!SL�+���C�LKI=�e�4����6�\�^t4�c,K*�����ؼ�%��a,bކm��p��ܾ�i��La6ܽ��,��]A���_\K��9W��M�T������|Y*����1y1�MN $md�F��Q쾀ꨄ4�o*����<O��	��mZ�b4��wsC�KQ�ۑ�_���_� ³��E�P�Nv�5�eu_�Dcv��T� �!��=��,�2u/ق��$�*�M� ��S�˨�q�_�ׇ�73������
*T�g�qXx���h���3�v�3֝Fh���!1 �M����w,�]v��hJ��v;и�J�UH�V�x)����Q�����w��,�?�S����vПʺx"��C&�����c��]�?�4�
�x��҃/p	���b�Ą���8LF�񞀷L���ʽZ�C�<�̬f|�J|D9N�X��G������_�����}_ͯ��b��4���$.��<�M(�ǞF�,Lcvʳ�k�����:^�pDoS�ϠN�$jǻY�_��,��%!Fh@����n��R�9�T�T�U�M��q1i���a���a�"`h�d�Q�۬�d�����p:�}���)�Z�µ��Y
�kR�V�����@t_�,��_��kZ����}��e2Y'�e`������,WF]�'9��=��e~��o��#vM����zP9j�*���/�cIO1(�4P)�6q�N<��t��E�����D����U�^U�����~�~6�����E{p˳��㤺d���W��ߪ�g`���ǀ�V�(
�|�f����A�Cl���*p��w�EF��HL�J㎡���n=p[��b3��t�!8�G����$��	�E�Y����
7>.��\� ��m�5>6$�.��Y����,6\Ƚv[��0Z�S~k p�N���g����ef�6�3�I��R�X[Ǖ�Y��W/�ײͷ���mь� ���^s�C��t,Ɔ����޼��bUߣ �m��>��=R�{؝Ԝ�(�Æ�_#AhRЕ���FH���
���]s��t���q���9K�c--��и�E��L=���"w����ħd�$i[q����P�'b�p���B��ͭ�T�<���._��+�=M7G��8$��/�*��%�+!���./s/�3�~�V]�x��=í�v4"L�F "���a�S��`:E~L�*YH�QN�?�I�+L�{o�-�T�҃SA�v������Iku\0��[;��+��2�E���W�sI,���21�1aB��(�����߿�t��c��yR���ݕF�����6Y���<��[.�ot`K��>A����L!��.a-��vv�;Fv���I�ZM�̂$�����?�k£>M�0ıLD��wQ5�v
 Z�0�h���.�����1�(�6��U7:�iã24�~�u���4ۮ���k}�-b9�e�Yp} 8�rJ��U[[�^a��h�lz\�f7�#mbF��]��<���V��u����{zc⽵�{\��J�B@J��_a���J9�B,��>�jKM�(���-�X:ުI&�:�a�~=\0�� '[�Y�Y����.��`㈵����0j�%��W��#3�����q8V%����E��e+���F�s�/&F�G<D�a_���& o������v�e2���ip���V��M�_���1�����~*�y]�E��j/3���еȻe@��ڻ((=�b�|�c8��w,�y�	��Ɏ b�n���L�`>�H+����)���݃
 ��,����xH�v�H��Q�,����`�{�ɺ⍽tUNۀ�W�&"+�V�4��Qp��hRR��a��)�?��&	�-���Ȳ5�	_>�,��K����%8]��K���UD�4��}�_b���2Ϣ�aFo*_ܥ;����$|��Ơ�9ㇼ��1.,+�h0���~�G�~GMH�C���}�Ȣ�SY���b��$q�|q.c��g$>�w�*�'�Թk��R����G�n9��f����G����s�{-��U�f%0_������x߽%p�ժ���������F#�0PG<�@��Z�2+<�4Ӊ�$�k����L�[{'��s]�(u���ᨋW�!	d��.K�Ė��]I�q�Z|���6�����(�ΠL�h��P��V�-u���=tX~�-���ezq�j-|�49a&�d�5�U���	�f���W�H�?����X�,����X�?�~���͑�(ߎE[Y�� ����C�sXٳ���'�=�%
vW�i�2�<`�k!LAıv�ѻRJD���_QKw}��Fd��]�~�2�#	���E���-����`�'�������ީ��<FT�Qӣ�������0GR" ����w��Ή٪%\��h���v���I��?�w[/ 5�q����e��W����"���lx���I���(d�$]�����Ŵ�x�Kca�V�V�|��
�+�f�������LZ$org`�y�c�|7�1�3��r:]8�Ϯ��9��1����G�k�A�[66)�tSɆA=�n�v��W�����s3�b�a`���I�U�P�<X��%K�Jr(E��}/��!r�����5��ϐ$<f�	��w��_B%#��ɚq�&C�s8˃i�e��Y��@̣EZI�/(�eĆ̳k�����w��!C?�Sv'�q��Cx���U\#pA��b�1<2��e�L�PȘqZp��le����LW�N-Li�} *�Se��f���$���a[!)��E�Oy����ĸw��/߱e��P�f�����%��G���Μ�N��#�����t�ta��S�PY�Ѿr�&Z'�s#�.S�.����d��^�[Nxמ���R'�X�%�rڼ�r��a�"s#����	g���^p��غ����A�6���aGq�ǽ'(y����2����Bœ����`�����vqYn3lPP~��1ӎ\�+}u����A�U��őC�ݸ�����Woq��J ���_#9l>%F��פ�v����������>�9{��cOv�����c��uwI]�+]���Zm�Y(��5�0����LW�����N����PU�����KȭI�q��a`�ׂT�_DWI�b�0���͔�,��(��-v#�hO�����M�E��DKă���O*�f�(��_����x�R%��Z:�|p]�zv��$�lչ����k$�^�_�J���uNWNy�Q������)$�7�'t)�1�f��h{#k(}k�?���M�[s�~^�P�0����0v�U�VP�O����\������9��F�š�LXL'>��XNC�mrJmC�Q	�
�L��5; �����P��`���D��q��(�K�'럘"�y��QcX�]$; ��|��@ʽ�������J��b���(_%�֗��ײ����+��
և����a���Z{��50!�ޏ��wr.-�{.]I�4�~��ZE~Fq~WBQ�����+��תs^���xf�s�rV�at����~	�ߏo��;��ҡ2��Ս�L 
X\i�i#�jܲ2��.�=��ѹI*��%5�\���[5�m���~Y�c��{g攖�����g�b��u<�B.�\>:�9I����`(�M4
�5tk���N��SA�+57��%���f��>
�H���ڷx&��������M!���*�ժ���mu'%X��U�C-ZDS�q�A���,��J���f���b����0n�H�":k�C��&�`����x���Ov�	�P��)���w^�Y�hR�f>�-f
�g"=��rEp(�I���ָ����7GY�[M;	W%�̑���G�;qs)������	��qQv�a�d���a�/���G��/`P}:���Q����) �m�H��om6����B�Ҕ�r�l�����]a���ܞ���B���^�9D�/�ɴb�!�pn�?�{^�K{4�t��?50���D��g�uS�� odI�Q\����h����A�_����^�GuZ>� ���3B���BQ�y�w2��;� ⣂Ԇ�K�#dEk��Ij����������M���Vep#:�6mJ���!mN���K�
ߊ���?�Z�X�M�X�w�^�YNۏ�(����l�O�h���5���+���|����y�X��,�t
:�:�����lԣ���[;@e[�>T��Ճ�!�*>��O�7:L/:��+q��F	��`�	��;�HQ��݃��u��MTU�>	7,�̺�޿���U���D4�uH��D(GB�df�TQ�����%���^ԑ�+(����/�,
xE�6�EkP�0�ɲEh�M�V����-�;�rq5L�G7[�����+i'h���7%�;����N9͡&3s���-��/�wC/��e�]&�PP6Ft�.���"�<��z�4_������X��T,�4$H���`�g��5����q�\�jR>5�����UIVE�?>��s7����`?3��\�pKL��y1��,��d�&���GD3RdI�t�ƣ�PujG�(���	�r�;d<tF�FMT�� %c�\/jx�r�/�B��������H�c����3�͜�~��7�&�寅:�)�S�g����uc�@����bŕɺu`��?f���<�)��BB;�t��=���4r��$��eq{�[��A	�~���2�?�����Wf�j��#AW��lܯ�ʂZ{��T��`oٙz�^���ԥt%�h�3��ծ��t�i�^�;y���z��B�z���a��&���[�$0�Ⱦ!\"W�K35Y>x�\��\ɟ��=:�] �5�|�2�wZa ��a��6҂W��x{�+��h�o��&I�<y������$��ռ��M��@k��y�=����=�
-DH.�K�&Z(��k���AB�Q2���\�AG��)�d��P��}s��fޟ�����o�o�^�y�x��:��hU>���2�j�\��A^J�4u��	�35z���8w�o;`��(�d��~d��G�P0��u���u��?X�rI������L��#�~��E�Ǐ�k��Ѣހ7v��e�M�]X�=�����Z���8�ne�Q]W��J��P� w0�Q�V��?h8Z]��)�~ܱ�-���(�@e丳�jёҡ�π��N�]f�[ˏz����Wno��\��
~��n���_bK�b�F�����)�9l���R�n�Y"�;N�@Ӿ��)������Qg�5Sn�?�q�3��/�'�bY�����nf�����o�\���{��ّ�դ�N�pn#���h��t?̵��X��\�I�H_B��A�ܭV<X12y�aU,�8^��#h�K���i��h7���l�
vk����������Z���{
���H��w4�BN�Z�/5��_�y��66l�>.B�K�&lV�DD�6*���*]�f��8Y�DU��'5 j�.�huR��	d4��)��տ�K�TZَ�M���SsH��O^,[�^y76�o�r3Dm��wNP{���h�o�0�����K����+�JV�.��Cpm��p���?�!&�B 5S�Ji�$M�3�3�����6�?6�R���L�{6��{���đ�g-e�iљ8j���5E�)Ѭ}&W�BB�$�{�2�@�����L�i+��CF���D�1з���R��ԄoLs�-yw�iD�w�c�K)��������?N���g(>�f;�S5 )w%B�*��� �����:��`Bȩ���n��ѻ����I���	4n��Wɸ)6Jp��_�^�F���qO�3@�Y��ih�1ŖH ��{謲:�_���'8u�8�IW���	�S����j�B�h����0���~�x�A1�����~���:�\ǖ\��L�;��+X���'�Ro�m�*��#�{o;:�VsT���W�Y���;�e��R1���6�^??�nZ�xs8t���M��@�Z�(�ON�I{����Go���NLa��$ ��HU��p�K�rV{�f�`!N����π�M /����5��4��֞V�3g�t6���W���y�X�0sdo��,P��#g\�ż����3.R���=�$����v�h�tG���-�^���DU��4�xʯ��D��R�Ď޹��z�PB�'�|���o��LfCX4-Md.�F�q����9�e��$��t��Kqܚ72xT-ဵ�s�!�dx��Z��� ��Ղ��ݠ��{�Rs�w�$_��I��C俢��F�ʞZ���O��Sސ��&旀$�G�N������|����H�i�9�9L�3�I�	�pt���
+��ك3K����:giT�]с*k[�*�G��� �],�x�Lk�3��x�1+_�4���*z��6U�u�@�±5L㲏s�zn��������K7�<ݶ�ɂ̘Eắ@�:Qt�^��<JP��>��$��C�����dcje�0��3��ľ��v�v6-���m{�4��lo�:h�^��/�"�V0t���e�"��и�p��Mu'��ՠcDQw �#TB�y�s�A�.��yd�-~�<?ב��^lN���mG�Q�b���ǺX��ߕ�t�`�ׁ��n!�I�U��0�"l��R���9`����v5ZM������wvkf�?CދB�p���-�h��e�zH��(/��_밈����;xΛ�^�j�l|�YG����H���.�ڲ,���|6���Fn�,ʿ��\ؐ@ا��;:ley�}�D#"l�l	�����=�w>�X��*D,D��[�@-�ж���*ݜ�1�]�Ռv _B�bC\�P�\8J�9S�({�+d�1�l�蚖Aڹ%������S��?2�[�v��-�{uPП�kYt)vυ�-���݈l�ܪ��9���J�I�,��a��Ƥ0��z �G0�2g�$U�����1�M���Љ/8�ŝ��p� ���"���;��{��_��T�pw[Mq����z��nT8]-�AnX����_�>��ҸG��q���+��~*������(Q�^ѕ,������	�f��y�5�Ԁ��@�#��!�$��L̝����xtc�$Ud�;3�@�>�0e|��&M����]���b�S�����(����3�h#l���zy��(����-���B����nď����!�������(�$k���aN �J��P'w5���B�����i6�[#�r�&mc뼆3�0���K���*���Trd$� �[t}�B��#:�wG˿���)�����QFP�+w�H��~����4����oV�.ۃ�&x��VA%��#}�uP#�%�XJ�8����"F;�\�[�׽�1�c�Ak�֤�1}��??Ù�֊�&ɼ
wL!�)�������A�� K�*`_�Y%��˯pqɛw���F͙�:���B�Ӝ6���~�
$V��Gј���Gh�cLN��I��(�r?Tӣܣ�la��q���y��?� ��ҙ��2��K/b!>фؤ�`-�A'��H����H)� �A�Ѓ����e��d��R��g,����ڭ�_��ν|�s�g��I�)�_���B[��~�}�c�=-[:nG�D ��xg�\s�ӏ�{*��r�����[�z�W��3���C��p���3�,~�d/��ncﬥ���e*�ٶ���g��D�2�KJm+�����ݵVB��r�L���T%�*�ņ;��A�U�;�iN2��-�V�.K-a�	�u�q_#�!��8|Ak.�05��J������AA������r7�^>�W}�ܜ��iB�Δ �Q���5W��A�V�c)Y�s1�W��J�����z搧0r��S*����w�E{�aά�A�� u]�u��PX ��d����f���}ڽ��he��;�����$YQb

wQ�Fb�mRj�@���P8�����t0��B���͠}!�h7�e��ĘP���� g�f
�$���+������`d��.Q�j�$� $���"EG���8���ֶt
�;i���TF_����\ߧ2�!�2;��/@K^���̒J튔ԁ��������߰a��7��n�T�s�6���g�T.%G��[&uY�[/v���y��E�e�<�3[7$��L�ԃ�Y�����p;�op<9�/��-=�.ml4�{.��i�k$>�*^��w$�2� �/s���j�{�7������agp|���; ��6b�<
�}��ʠ6l62��d}�d̸��������Z3��v��C��� q�O�s��� �o��ԯdpG|��za_�Mή�ce�EI��y��@��@h�ɏ���P*u�U��Іdf ���N/P�x|9�;N�[\تN����k�iFg���FL�pq�4]<c�L��k��}-H\I��o��,�Tա5IR��4 ��ym^�㷀A^��B�L��9��y��=��k�
�e N'�s;[z��B\Yj��xu��eVIj%��۫��(�U��a���zۭC�f��Ac�[�J�*[l�`�M̕�+���	O�͘�C�-���wfeG8��Ѿ�<]OEH��۬�ێ	t��D
`��.J��R+]��i(���(�^�T��8r�� u�cã����BOQI<����W��
К@ބN��]��}'�^U��؉�W�����<�='v�cd�bep�b����8�%"��;N)8�Y [���Y�3��zݱ�>����hBVɸ��b���WҴ���P�;ج����Ծ�~m �$O<�y�\�y�/.�����S띝��$$�M4�x���]��F<�#�g��3�8�>��og���ţ��lq�7U���|�sf�HZ5�ӣ9�^=9�a�R�o��e�K��0O��ه����\ z��~�T}�d4��w��si��m}�)(y:j���X�.����$z:?�-)u�)$��'���MM�߭��Pm*��w�����-�~�*w4�z9 MyQ ���n>���������=�Q��S�&�q���h��K�d�d3<��YN4������8���z֖GtYl0\��wg�g�<`�hS�%s�P�)A�q(�nc�5�TLļM͊a���=��_F7��u3r�W����`�W<�;a�����ōctn�ͼ�u*�	e$U0-<jJ��A�����L���*��/H~�*y�)�ʜ)\'��%V�N3\��n��).�6�6=���	� �=Ia7�bA�'1�Ek��l�T�>�����i&B��_�s`�a!� <'z���"��,���+�;���
a�.�f��	i0EOfpw?��i�n�z�S<������,«a>�xލB��h�C7��ڍ�)�g�︡��|Y�6S�I���?�G �x���EFS,�����]��1���q�f$��#��i4b~�([L���=`3����NJ.�}.��"I$���r�g��@� �4���'��Id3�xs>���{ENﯡ*��69����%��wh�V��ԅ�~��'w�%ݸg3 ��/̢zv���qS�|��8<�*1�|���]�h*Jg�vQ ��-MyG
�����+��Ll�>��{n2QD
�7'D��CC�b�WxU�s�3w��.��R����c�C.����W4"W����^Bh�_�|H�9�o����c���bݟP�_�Dt��mR�c��g�
��|̰�lt�$y��� �`�pL��� �f�M�л��e�-\�?��a�P�8N����Pp���OHwQ�U��(�)2�&�k)�~�� �P��A���������NAM��D��ߪ�W�>r��۸Ȧ�����j|�ى�&�V��pqٳ�_�(�;G����u��N.��Kt�����{g�?еD�dE�p�(up��j���#D2���C�)@�A4t�[�hD~��Un=Nv���ʯ�~d�����@v,+ N�pEG����Ho���P@�������lЉ���@���&�U?KLǚ�Z~��ӛa��c��o�:7�ӈ�i�����%%�B��C�����	��x&����97pr�� �����ٰ��q�b��!c��4�u�(����̵�>��.�2l�)Ƿ��d>��7�o�q���q�O!� ,��bi�@��2� ZZ������T�^�cTxT�28�$/ky�3�ƫDI��`?�v@=:��9Fvo�������?e)�K�������k�&�[3	@[6:�~^4v�~��FP�bC�6L��k-���]@yX<�P{��Ain���,Z��P�F���p�S>���3�]�ҨPs�Bw��%�@����F]*�$R��6
:Ɉd^A����ҹ��6
��4�m�
��"�)�WV��P85$������t��Z�|�  u�Qe��xjY�c�Zs�9Bk�\N��5L�/�Ӌ���	(�J����aL��-<L�m.�^v*2������!��œ�٢&�s@	�v��J��ˇ�*�Ο(4���飶��!�4EM,��B~O�v��}����o��8�ܙڦ���"��q$���z�R��E���&��ٯ2�&���C�l?�SP��ڪ�41��e��c�y��x@+c(�?�O�u!�6�P̌˸i������s�/�4��(�� �
k�����FC���9uV]�6=vH*T�+3W��fL�N	"���|H�NAQ����˷u�X�Y,�`�$
� �����M�ٟW�28Z\h��~��Q-�1��Y/!9i��ZN������k݉І�f�5ঢ়��	k�~ɛ!.)�xj�U�$�m���Bk��Hp#�Q�~b"�$����Z���Fu�#���drҮ���͒Z��u���}"��(r�t�̸��`� �K�[���b�ad�c��a�%�]]�v�0Xmۙ_��=e�/FF�<n�L5)6F���Y�C�h�@���ZZ2�V���~���.qM��