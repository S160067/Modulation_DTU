��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����>�S��fI#�l7x%���$or�#�6�y���N�i� �D��f(�:eǊ�` ��S���^�mBƱYjA���v�0��kh������#�v�(#W��ux��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>:��cG���Up�Y^����˚;���"J��+��sc��Y6�f$6�5&���z���������`dcR�+��b\�v���D���ղ:h�W��j����='�5Cq����7�r!��:l�6�Fo���_˪��k��LH�]!��0��W>^�f�2u��uu~�
��.��%_�|h=*�����T�PB;
!��ϛ�����cQU���^3�kM��i�X�:)Ė�p�]��tF%�/��P��8�+�ާ�x�8����O�����2�L�%:H��nIg�XRr�a{j�D�	���<�4T(a[�WzRY�&��)[���V�6r���e�G�|�в[��H��e^��2<���6�띀Oz�z��d��R��]>�֠��BZ�>��͍�v���yN؇k�a+D*c�A7�euBֶ�v�T�� ������D���|��ʥ-�6��i�m Bӟ�u�=r�h��L�V��Yw���%X�^��X�{�g�j��dh��/m�7'�ď~U�������� $�$��+!�� �<���5�����kǸ��)�����F���4��i�ڄ���Zpb�,|�$&D9t~:8����������hk�F22;�}�V�/}�F�:H��n�<4I���L�.i�/�z��Y�Pl����8snYP�o!�-ɻ9'��(�[����f`uA�P�?7��w1���A�`:���Qdr�b���V��KXƸ�ޛ:�?�drJc��ďF�xF��l�e���oI��%./�c��QZp��߹9r��9�p
�3[�J#yn�Ϣ�[�V�dn�����}�mo-�{�h�6��_90�iE���0��XF��%4����k�@�N4�ᅦ-�R�_����a��ė��
w �4[��K���e�x�Û�N(Eo�SX �y��[q+�*���]���ڣ����2�L_��;�K�1�qN$1���s*�_CX��9&vm�q������{�-�$��"�G�NQJ�D�HB�Vrwԛ�Qp?��?^�2[[��(�X(�qgEH�n����lj���� ۹�j�zHqg,Zr�>�~b,�=�P��x�#k��|�j�����si.Ó�/���G���zPҡ�FM����.)7�	k A�X�1��Nb�$�s��s���ǚHd�����}�4p���a���eJ��S�a���M�,{SrXcw¥&�Ɉ����@$���3�Z�� �(!1���BHU����y����\q�=�'��:��.EG�S㾯�tѺ��=�)CO���7���hvV�:�MRJ]��?�/\��P��$��yK8��3�5��̆�ǽ��W ��x����+8����:��_��m�+��N��(o�z�2WtÍ�3�S�zV���yz���T�-ա���B09�_ش�YD��|72���S�N�Uj�o���/{��R>֓F�ϖͶ�
�T�8D���1�IG:��T�&%H����2̧��l�?��q�&z-������<�I�oG�}	�����6���K���C��QX�`H����+�#e�䬪��g���|`�3� �m^�0�<��Sm�oM��f�!��i��Ыv���J��8l4:�SGD;�E&���[v?�b�.&�6!�ġ����
��3^�� cQi��!�JJ�㎣͍�6p�c���(�ӎ1�]r+p��-ǸW��\3a(�R��.���L�7�\T?[l��<�F���v�Xp<��;r�tv,.r/��b2�6`_pU�i9^���ə!�4�uj�2�Ǖ'��|a��rK��ŭϸ���΁/{�O	�m���0��
���sr�k��?��w����*1�*�q�
� �h=
O)gfȎ>�ܤu5�t� �եɛ��	/�7���%)��s<���{��53��<xh9� ���\cyn��h��_�1��<.�Lr)<��<�?]v�NY%ӎ���T%�L�����\-r�J�rߨ9�q�D<�34e/�ԇw]�
}�s%�||}iͩ���)9�p͞�f�)=[7�*�R������(&ޜ���'�6o�:���;j1HJm��%)�/������3��0����י�Y��hm�B���7��������C���e$i��^z�"1��h�4D�M�˕\{�7�8B4��G�Q�U	��ܽ x������>D��6A��
�"�)�>��_lM {��&I��_H��¸mȳ4�X���e?�8�/��gb?$��X;��z�!�{�)�k�쮙�<���b�b����ݣ�销����^�F�|E��iӇ��x�G��rn��:́�`o�������a�e�9���`;�;����1 �ƾa;ͪh�	���-�cMl�[��B���F�c��"&g��'�y��)|L+��vo�;g|������ui��9�#VY.�����~��n������i���!�YD���D?.Jg�����|�Y��ħ�nX(B��d���'�	�A��8��Ε8��-��eJf���H�\�y�c#?�Jv幇d��}�7��D��������@�@R��CF	 s��b^��#5�����^���l���:k_�:.7�j|��}*�3��v�����rں�����2:\��tFx��/
*]�Zp��8U�X�����&9ʄ�����-\��tkwQ>�k���xj��I�@�O�y�▣k�S������o�k�6u�\8⺮d�6c�B�u��@s��j6�#�g}O����LM���qж�V�Z~?{ha�@} b�֦KV�:ҝ�_����L�=�:_��@q���ru��,����b\�&�:�6R�&��a�_U3>�»)d�v>�y��\���o%�?�A��Q�"�'U�l�0���<^������+K���%{+d�h�\��W�EA��Ӳ��@>��V���c��������O�a��W��m �a�KU@",ft���h�tU47 
z!�Y�<n`�)���,�B�NFZBY]fI�D���򵠟h��D�{�\jT�^&��5��@�VaM\�A<�}�hAo���H��(�׽?^u�U�0�q�Љ�x��.����}V�d�Wfi�Y�����C�x��9�vx��.h �I���u��n`gs݄U>�9���D9aLT���ގ=���ht�c�d�:2[v#��]P�S�#�
u��$T�� Qg��h.���� ҁ��ܒDMOlh���!�=�R]�kL+��RY��^�1)�6�.�6� E��;"�P];��7Ŷ��E@�&˝�4@/쾾��f�j�|d	��<I��e��,�Y	�Đ�P�(�3t����t��T�w�5>�.vՍrU4�{����2�.�~�]N%����T3�W��b�Պ�!@����V�#x+�#�;~"b|$��tF2 ��&�k�mj<��֧�?O�%���1��j�QT&Ty�9O��;�5e���$������H�)�&O�L�X�T���F(��f_�d��8WO�ҷ��)*F
��UC9�V����S���|f)f��½4���hK<�v��	 τ��P)e�X)�s�X/\�_�Am�B٩;y08�퀪z8|�E��Zy��d��&�5<TZ�4������o�CX��5�䂸?!�b/(L��~5�XRn�F���t��r����Yj0��m:A����bOry�{_�&�x��8J��K��*���0�*���P`+E7��A��_��]��º�
�~�5�q�h�7w.�9�>��Q�etߥ��@�H�='j9�Q�w]�� =�< ��6�3�� �����[�z��h��o)M�Ji�~ZhƱ;l�I�5=B��u��/�B�ʯ_,�q�dV�����Y1\pΎ�3�C��$8���3��Lt)_��5�@�a�F?~uP����[�_���D�V��kН�
D��[1;o�3��/�]f'WO��
�U!Ls#�K���籊Z8b������н!����y�����d��R�P�sPZ�c���F�eGl�k���\�0a��0���qi�����s�3�[&�,R�X'�M�J|����aɸ�)���2�$<�j2������14�V߰�l�ĳ�~1�)�G*si��Y�Xt���ĳCo��T�	��&�8�S͠*6��OǾ��P�$w�i�Jy$��?3�\3�{0�r��d�vG�)%*��s�����}�=�^�%�����=���H}�k� ��u�jYA8{t���QN��&[�2I0 � 4�!�]Vx6Q�{\��}���;�e3�g�o�oH�F�DQ�'�ub ��%�$T����o�T%ޤ���<�g��P0���2z�7�3���5�����	��{J�]�M23��Y��~��-���V5���at_#���=Ԙã-��Z�I�5�1���.�3����t��vc��4��M<J�z��}J����F?v�|)3�ڞC)JVwai��/�!o��(d{^���MY�ɊG�R)��N≍�Z�S�v�/��]�����pmކ!@F�=�3�����'wq�������fw���_�nw�i����F{��擠�R�]�����a�+�h��1U�͐}5�{LfSye���z6vuȎ,�Ytk�E�����7�=��O���C#�/K)u��#�`��H�-X�Ey��ؓf���9:�"���H��NRԇ$�a�8�!�2��AA��ݒ�_�k�2 ̑'X:e����fȨ�9��(W��,X������b�5F��^���^in���!B�����܊��G��&vAٱo�t�<gːq�ǥ�
˻k��E\�D֟��W��λ�b��k\Z4q?<kԵ�$�C��E��qzje��x��i�ʰ��˘�۲�
S!�����]}6�Y��Pt4�̹D�B�a��c�B�W�� �"ʊ�$>�)�z�T4�?I�$�;	)�.M0���ޒ�8����K��=$��*��I��+�f�����M�?>�->�i�̨C��[~s�o#��W��k��4rF�y�rEl1aI�b�]��_���[��4�b@#QO��8�R��iP�|�J
T����z2!��5�*gt��dZf��2��A�V�eȀ�Ln`���.��%�埞^�yY3�����5�my!$�N�:Y��Q�w�iK���S���੄ӇQ��q]}0��T^���~�����za���}��d��@������, �(�-���D��d�����E��r�0j��ի�͙C,*�X�R�CHp����� zp%�o��xbadQbuA����t� �����$0���k��a�]��e��7(�����@��+2�Ug�%*%�� %��}�e�	����<L��BW>��XF�&4�H~G�a��B4��Q�f�T�!f�y��4��ȸ���x��T��S��nO²M�1�ܨw(��^��7�O�l}��3�����Ӝ�<LȨ�`�=�ԊSP�=�+��6ĉ=��_��T* �^B�QP�Q�ảe��F��Ҹ�Chg/���F*�i��.#������
Xm���nlՉ�w��I���	�F����57��4�|̸p��t4]������T	�)�lo�Q�}�)�@�S�
J&i&��N���4���ʛG`�a���9tC~�	>�U��"��u��7z���T�����ڳ䂁�� �G�L���<�L�>�C�Cވ�N��3C�R������#j��D�|I��U�t��'�?ѝ2W�_��Xn�I�&��� ��[���1����-b���lJёc4pC��i�ް@�|[G<�IQ����2n{i�1A��E���;���Ο��CB�UάX��dCVsh�M"�2 ��LE��;��-ˣe�Z'Ha����CǺ��]b���Z=�\F���(�9��>���I:�|y�ok>Ҫ���ef��(@��B6�D�_Y�U�5��F������|g�	�AP4*Y4��',7~����-��\��=�7d�#+J�CVeu�F�HC�;�
����u�e#T���w�l�{(d�z����g}�2����tM�7���������FRB�ٯu8}��/�:+f�md�m�O��W���1�~%7�[�J}z����D�?fu�҄0������uA0�)��kw>A�>�f��_ ��/<�8��z�����M:���P	��1�!
�J8�+�Zv}���і�7�_��`BL�X@7�Y�����?��:���2|�O(�Y��!�]�r��d��sC���PW]WR��s4$�%��A{Ӑf��ad�o�SIy���M	�03U���߻s1���4��=M ?ji���r-,�^�����+�G��R�����`u/9^d�P��>