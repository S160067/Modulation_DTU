��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���,���`�Q �����6�͍	),�6�md|_��n�x�"u������K �5owJh�E��qڑI9����%,%UEwf�x����;.�9��p3��,/�֤����"��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
N�m�H2
��j�Y�? ]r��j�p�V�d�����띜�7���{o|��hg�EbVS����K(�k|@g���)��i���7�b���&nDo�/7���)�&	!%�Kw���qi����N�c����S��g\<�e(͕-�T�d�G�KD��P�j;��|#r����l�|�ݾ�SQ�w�v���|d��2�ښ����g�Ti:f�G�Ǐv��3O�o�d��*J=�#��IX\�T������2)�En���3h,8�Cg�-T���9�αI�4;k���N�� T�"u���P�aT3��4���F��x��r�gav�m� �ᡟϴ�^u)].i[ݤ���*�X{���db�#h�ϟ�j���(&>����,���1=�<�-�����ơ/2A�_ o½���Egi͡8�Ss/�S���5p��A�H��)�U� �aI�Y���C��u�Z��j��-��19���r��WbJV�������1��h
W:��u�a-г���D^p�V���l�U�n~h���ĩX�ӿ�o|�� �J]�d_O��V���G�>�!v�}��b*����?P_먔o��e���a=�d�C�r��&u�'m'�Vi!21��h��|~���Gk{l�?h{ۀ���*`X��E���q\� l���)� ;��c���߷(��q
�cl2"f�t������'�ɒ���+�3��;�����-���2���a��4S^�w�)rm����>�C��(�O�nV����ww���͕��ˀ+�WqT��
P�6FT	��V�����5����	�wK�9/��'��_��?_ra\d�ll<s�5��8�ɳ�4.	�PO[u����z$���F-�����ٝ�eBc�g1�=�E/��i�Q����asO�=w�׻�.F��F�^k�pk� �ք�?'�v��K_\n'b�u 4�G�oגџ��J�����\^\����F֕��iJ��͜6�Ҭ��0��EІ%$m8��3�o�����[/O,S�D���
�z
$��#���sK%�\���7y� �
ڽ�u[�V�<0�؎�Y�W��N�����9�d�̳��t [W�����
�3�K��Ð��� �Iތ0�F�xs�γ��u�?2�{؄���Ě9(�D"��i���3^�y\�H֣˳�'�I��h]��=���S+TBM�al�m��BR��8(t�	uM�4mYڶ%����I�@��hG�ϣ˩qG��邼U3�X�lp)�E��l7}es?��U�%(!Ϋ!������{C�z^�s)9�"P ��:�"��aH�ڶ0�R�e�c�mP�P�� g�'wt�u�6]�
��ԒZNӅ$bĥbe��I�A�Sʆ0�w݅'t�C�L�ِZZ.�l5���]�ؑ;�uB�z߽"@fE�*V%��dc)T� �*��fj����)�I��o�Q�W��+�^4؋%����*��Yo`�ﱀ��t��a�nΑ`�r�@���b	w��Y��j�d��C�D,��EH�| �U�Ѩ��SI_tIe�-�K�.<^}�]�>$�W��oK��(�Ώ��:�Pi煒p4w� ��ey���^��|H�L8a�v=�Б�[�a)���*��<�:J���9_>Z,���f�D�>�]yeuf�΂k����7'���TQl�
�=^�.#�l)H�4�CK��0�� �c� @���hEG2��p{%��E�U����Qw$&Y25�~��CsU0������Ӏ�SɃ&SL��E֔��ff�R ��q��9VEzn�z���B���{i��C`�$�����t�I���`�ȝn�T���+����>K��z߻=zHzޑr�h��q��T��/�wf���Я��}`;�(��#TZT��{���������<��*��fXs�j�����V�ގ�J�"���XK0�s��zB����od�i��U��i����g�H��4П@Ll>@��$����.B�W� ��R��{�dܕ�Z"�`l:�siCX~<�l�'6\(�3�:͓%�}�e=�s�CM5jbYA2g��ͽg���y2��FJ@��o�xb�ԟp�jMױA���(��L�<%T4p�3z>���Qد�����f̖ӻW��~5�#&)��������-c��=$�~�J!gh��y��"X2�i��v:9H��*8,F��� ���){��/@�v�-�ttX���~F'n�s�@������7�37��>ºɗ�����}K��9�Q�g���)G� U暇�(��(�����G�/�Y��A�7E�9��~~;�#T��T찕q�J���5QG��9g}h��гK�����<�BWhI��1Ӌ��dJKʕ��:�WC��1v:�l�J��V��/�mMD�H%�tmi�=0-S �������3
`�(U�ہDL�aY ZVQ��\���Ֆ�	��ER3Fi���1�?%�S� .��,��bin�c]��{�5��l�J9�h�sˋ��h�Ag�Ђ�/��&2���lfp��8K�;c�-���B���	��댢lyƱ6���	�����L�a�A�fF�Y��V��C�7xx2�`u��Kb��[е�5���Fs�ީ�1�~����ufWMy�cd$�_7�.QV�r\���ҽc�J���ū����,V��U�0	3&��m�|(}���&�X����J�?j��,$��q�ى?T�$4�C+F*�_m��:�:�>в�2��,�`�88�<���މ�Y��k,��m"�E���� �>� �c�f�>A�v��k1�+K�7ϖ*n����A�g��T�d��IK�J�%r���7�
�z���D*�JdbÂj�n�Q�)'��W����>��`���Y]:^V����qB�/r���ˇ�|���$;ō�*3�j]�q�L��)l���T�l�E�D�a����-h,fxW�\�6_�����t�k�T's>��Sf��'p����e��%�R�P<Z/u�n�<��F4/	�$k�*�M(=��W��WҘFcos��c)��QԛSoR�}�G+�Ĕ��\~7fg�qFO��V<@�M1Ez}i�`�k����{XEG�
���00�fyḌr�V�Y�Y�O��iLi�o�*A,��j�B�9��'�t�!X�^�x�����Dk���u��Oj�+�Y���x`#���ޢ�f�5!\��\�j���K�֜�/�=*�B�P���>�+�ѽḂ��Q����Ty!��]K���-��.-��m���V�d�**��ط7Z�u��>�=B Z��Z��Z�S�.����.��9{�q�VhB�v�v/�q�C�w���e>��^��L���V3D�dH�4�<cFA�Ā��2�����#9��!60u�9����w���G�l��ˁ���A�p�mS����yp,���V��ϐM��u��A�?�+g��Ǻ+��4��3��l)�֎o���[�� �u�B%��>m�<�\��7��X�?Fѳ��n��3����"��a���T�H~@m�A�ŗ��[�4��(dH�������A����!Z����"5V-�I��Z�]r�{��Ɛ�3}v*�<���c�qZ?��Q����E��n�b���M�����-W����Ð�4̹�V�E��!�ْu	tz�^js1���`us�qE½�ʫ����j�Q�����
��5��NF�#�=��#n�5����:��(�Ե�;���~Q�c�t."_�K�l��nI3��j�����R������yk�?�o��.����kJç�P��U�Z�)���c����e���pM3���v��jy��{<_�'�G�|�E����g��e��`A�HMy��hm�'��E�0����F�D�������6-�Dn;]4�O��������d/���>�9�A����s#����}�z]���_3���l�j��U��#�(���^|a�Nt��*o�B�U�,�
,m�����՗�w6M-�^f�`f��t3W���Nwtx�D����Z���q<�8H(��;��+����������f�;�M4����e�6E���@��y`U��H3Z�����fL����3�d������d)Po��kqD�a
������vk������+��ڈa�z�%��p�z����wqVo�)�g������p⮳լw�*������W��+�^M�O}��\����jH�2��	(G������wWOw]�U�Fh6D�h��<�FNrmA���������\eB�
��<K�qG�g���t�fyp� .,�e��ݶ�� /օ��#���!6�v溪+�i֚�B1�c��4v�m��%�\�[��(Q���X�=�~=��+ۓ��Z����]�W8�=��ﮱ���'a�r&�<@���(��1կ��Y�����.d
�GƳXJ�p�ȝ�?�9�vuU�`�eV�i�MW���l�w�#���3I4O^cR���3e)î�<P��3ȍ���$»ٞ�� �-OSfX�����)S��=��i�#�ja:j�x�i��.�~�>��:
l=*UP� ����:"�s�n��W6q4M}{y��Zn
K�:��A�U����Ԓ	���J�
oy�એL�%�<(�� *kɩ�Ma��/����b�i'�c�sY�dZ����DQ��{_���)�e[9��[l�ɸI�	�w";l3�_g}Y�� #�ڧO��K;�u�"qXBx�itoW+��u4p�/����N�ywR�����a���v��R�ʙ$0��!���>^IW���ƽ	���[��ad�ܾ�p�w*lC���1�a�&� �-����n�'�yԀ�"�䡕3�3ӼؼF7i�f��v��+`U��@��=$�9��Kۍg88@���\�G�<,�b[b�,u��9G,k���
���%�'���<$/]�v��7�H�y�62V�����<��\B�&L�$rn0����_2E�s��-�0����uW����Bm�>+^�=���k=�1X0��r-���t��;�#B�)��x�������R��N�Τɽ1hI�s�4/�dY:�(�q����&o���&fF�`�DPJX��rq?v0��w3�k�<��R�s��I�K$#�����y�g��1�yvwDêƈ�+�^�܅�*?��@��%�gv�	:2��e^�]��r�����}_������^�ʪ^6��-���v�z�+z3��=��T�\��~����&��!�]�����ebHz��S�(��<%7�)A�da�e;�R��ӎA�����@����HYe�X�L��?�Ĥ�����<�����-������z[u�J*��ofЍ������	e�oy�����x�L'�"���L/,.��o�6�{��'��*n�o1fȅDm�z$Kc���1x�TU���:�L>�Ưȃ�F91��LP$�_[ �u"|��Y����QS	�Mr!Λ9'En&VR��Y5�	O��x��q�������o?���R�v�j0y�ۥ!<��s��*[MX͊�=A�O���-z��݃R�ʚ�������e����$?$���i�N6p��D�2^��lc��Vj`'�l?e��缴?�qpS���)�"ڦ�y�Ҙ�;UG\(�9�2�Q�LC��~f�C1s����{ �yfٰa�V$/���E�0	:����yZ��*�$��Nߙ�!�ω���_I�������n�FL4v�I��hl��J���a�ao� Xf,��I����&�@t6y�#�Y��z������$��[�z_@���쉪���V���,Q��P���J'��W�׃�F�-�����O3dE ٌ���r�=��.�/z���}�.�ߢ&����g����7��L?�u{S_�:h?iJBj�<�ܫV�H	��@��W����b^ ���o'�vr�V�?,Ԛvg�I�:[�sD��k'7ӚW��1�UO�Cl;��L{�Y�2�:H.�`N�);��3���u��<}�vhaԯ#�Z���m���[�y�6���~]|q���k����2z:�y���!�x%�7o�eE�Ղ|�w5k)�]94k_�`c�uY�ܖ���H��Hu��N��Q!+�z:-ӹ�JT�`����m���C׋�}�ߜ�^�D��1O���9(>���Ka,�qO�$C��%�]ռֹz&,�tH�hl��1O`�, -����0��`���v$G];��� �]29W�MGuҖ�d�C:H�+!�kQ�ϴxt����4�&�yS���=Q�i�(>��P[ȫ�������&�/�`.Ӳ��ps��#����2!�H`Ɵ.�B~�\��t�B�}M�xd��O��JK�;�i+�L�F��a6�({����O<��ae]��CP`ׇ���(5�ڴ����sq {y�1�<�)>��Z��ة�M�Au 	90����� �o�Ӳ��.�WA�ppDA4
�[�~d�멘Y)��,�������D�{����ȌHp;�H{���T6Cn��:(!c�g��eu���g��JQ��^��v�-w����Ӵk�%���ڀ3m'�U(vF�*Q�d-:§K�=��ʥnFF�q�[�=&#k��9]��߃�� @N^*�^D��U0�Effo��������^�L�bȥb5����J���v1�7�c����Ե���;�	k�<P��9I�5�9�����Q�g�|6�G�Դ���=��{X���8�AE?|�G�$��*$�7}�~��.<�{�z`b���4�'��V�L�Z��(]v��/�gV�BV[o1���3��c�w�mE��l�����>�z/x�7l���V2-$s���p� �WڙJK�~>�t�+��%gcN� �����)j8z�;� L>(�í;Nc�9�'<�m���Z�PCX�>�q�&Î�+WÑ�������1Yd��mM�)\YR�_�"Z�4 �Cv��׉��6�#
\�vS��˽�-���҅��u勓�9��G|A�F��P��Mؒ)�����IS/ɔ�w����J��X��Te���;{�u�f��)�z4V_��(�Q��X�8S������7TF]�מ*�'ܛ��X����H�k�Gx�@@��ˀ��lu�"R�,�ک�v1Ry�������4���		G��q6���GRw���^wW/��FX����������z�记=s��FV��C���s�����G���=�%H�cd�?mmQ�+����7�>��B�s��WH����&!�T�p�B�2ʧh�}w�R~�}�0�K�GřJ*Z'i5��
�@�-���7��Q��TۅK�ߗ����a^�	�gGv�(�u��2��]f9�s	M��}R��NO�]���?������S��j�M�υ���*�+��C��,<����l@��e���li�c�	�s��Y��%�����7���K��'T2��ɞQE�R�}��b*�v+$G�6Z�y�]��佧��&�Â�0���qԖKa���l儓&�^�Q`#��2�)/��J�A+b����\�����#�Y�Q�+4 �t��GL��y��9�,�B�B�L���>�����2�#��D��d��P�"$>N4w�I�����R�����������t���Zg=]��f�V=���������_=�o�6�;2%�2���Z�'U��G�H�,�6��a
���s��� �Qb�v����w���� �:U,�X�ga�i!���5W��+��?�H~�b�9���r;�z��KT�yd�/��Af�_�?!��w.��z��.[�b��F��<: yy,�i,��v��������L�7���{��b����yEZJ:��v�����~Lף��8��$ �յQR�r�w��Yx�XF�����~��C��e�L�Q�A]�~&64���^���zC�)����n��U��El�؆+BuJL��|JTF+L���;dt�ɂ�1f�x�ɨ�0�B��̎�슏L�fXu�;����Jl�,t�Z��g�6$�
27ˋBaN��;�G��q;�"N�Q����f7&~c�+$�z��q�f{�/��w&g���K
<�1.��k�,~�Y	)B���RTT��
(��vUC��gNw��<i�fl�.q���H����p�0�R��5t�D����:�r�1N���s�����tč�w��s*�J����20x��&84Y��rԑM�䮹cu�$���G��,+��3DcQ��bI�ɛ�!~���C@�e�MM*-|�囚p�_ ����yvU����z��3�z4���ܵm��@۶�&t)�b!�b��! 4��?�������?R��'�>��ԧ�ӪS�ֵ�_+V�����W,Eǃ�\�֭� �[|�yw��u�҄c�̓�`~,]�$�P��jްuEϗG�H�I�۹�Mr�Qg/9{=$�ul7p)���&�F�$k	��2�[��7��|�n;I�w��_����̩��he_�u�h(zEJiHJČx�Jω�����2V��J[�]�o�r���\)��)�y�;�.�Xq�n�.e�GYW9�5]^"�)��&�������ᮋΤ���S��5�tH{ݲ[qL�%6=/�
���4&�I �x������-8#�Q��*�~<�C} ��{ת��Ne'g[�AXV�N�_G�Gd��Bt��n��Eڃ�<E�PaUӯWˉ0�#Cbx[%��Q�_Z��ؿ�a�T��:�n�6w»��_}z3+��qV윬�vʃ���k����k�+�v:n�b�.�~�,ܶ�#f�1$�JS���W�v�џZ�<̊m���;�UI�lv�%���xZ�|���_���	Vv����� ��r=�s�2��TK,'�Ƨ�ea���2�k��RPjs�a�30h5�Sg��|ffl%oW)�{i5�g��A'��<0��j�����+��P���"�N������Fx	4h2�' (N;���Q�zp!&䖖 OJPI�A
ؐ�KU����Z/%��`�Ύ�g�.~�~=�	���jP���
($�X�"�z�3��ݯ��_;R��`y���&E�!&.���ב��
Ӌp
lA��)�Y����Bہbh?�+'Y��S��MiA"��� ̞w�EU�/Y�԰��RK��ߞ�%������_�~Q]G��2N�Cd��P�;*�˿��˥γ�E��ժ�RS�M;��#�KnR�5�t�G]�5�c�
��s��4��V����oSc�|R`�y���,����Dv7I�(��9]�k�L���K�y(�L��׬_�A3�Y�A+���Kύ��;��ct��V�ܿ6�����d�׏#�y� �/䯯�T��h����(n i%Ѯ��c�Sv���Y��K瓤.S��o��=�r�3�Y��2*tL8)�.���,y(ۜ��|�ҍT?B�[,�'�|$�.��3�3C�&Vb��u������'�k���5&����2.gQ�؂��LH`��-�[?�,.�����v[��ɟvx���83<"�FC��I�v;v��2����O��Z]�v'�)L�r���ч�%�
�r�8Z���bsw?�_K�
t��k�����]P�ɾu	���� �%4g>��]fd.0�.������)T9��H��|�vr(&x�&۱�A���G5��7lt�$�{5�`�`l�r�R�-#*h?ɑ@����cÅ�bi��z��
�a���i�V�~X4�-��ėl�߭����ߜ�%��8��k�d�آ��f�E�D}lf����fxe�s��y%3�3�x���rZZ ���m��%�w���#g���>�\��$����������OrI@�Ӟaz";�<���;��¬j�1>Z|<�-�9����󾥮�hYMH���beL|�BN5��H�5���F���3tN].���P�o��ų(0MWd��l��EKV������]����k�V퐖o�h�OO�y�i �R�����%Ҋ�lr�/�Q_���ºXJ�77;��ƶ�N]�a Mp`��W���]�=c&�CR���YE��r�/�����b�n�?u͍���w1J��a㱟��@�p����%��n^�T���[����E�tf0�6*S�e�Bkz�tLQ_u�zvO�f�|w���j�.(�2����{�2��9^A���ί+Te&���"8-i�?P� ��{�O�%�|�""mTzwj���FS�^������v���5d�k�M(�e� `G(��N����1֡/Eq����wH���}�D*�Lq�.ML�@�������=�3a��R%�$f�S6//�%	��>/�4��C�񋋭����.Z_;�p(�쭛��Up���J'�Ⱦ4�_����ѵ6�lp�(v�,F���BD&�h?�"A��,���N�FPj�������םw�-�-��Π_#�x3��~}|1�F߬��6%���g�RT%/N��5��.��O(I� ��t^��LsVB�;Sax�F����ԂOs��<�q-cb���K�c�	�;-Y�E
}{���-�>[ ���cY�!�+n����{�T[���k�`
�@�]V�]����۲QH�{G1Q5~������]��Q�-��ȓ�W�e�,$Te�_^����>g=2Z&����I��#}��7Ѷ�l*�M����a��&A
���"L�HF�8E��7=~�l���-A&���fR�p!_�&�uR������1\/��0_�~:B�vc�2�|�/?R�n��}4W[���y�2. t��K�:%!��TR��4+Ѹ����W�!�����&_���I��^��������|h�I�,c�p�B�����Tb*,&��Q����V	��{u�zĸ)���Usd��WG��צ#�.��m"�0G<��d3^*N���Zv�AY�6z���8����sO3��L������d&�l�3�O��r5��c�9�F\ڧ�����=��%6j4)�*�Sp5�[ �Nc��]p�~��!��q�c���ۨn<S�$k��`�f�-t�˂�Ȗ|�SG�r�F��R�z'I10yu���Q�.�0YPC'i-ʉ�)�CU2=��+\=JvH,O��S|�|x��~�%E!c�4�����yqhtOշA�o"Н[��QY��yK�hX�W�,��(�j[`xVR���Q7�[%`�S=�nDvKo��/M[@�D�0M��L`
 �c���T|� �����������Bt�77SJ�ע&���pE�YhN������C��Z���֌����jbD͇_q0��B\(d�g�	�ag�������C�e���I�j׽�wP�m)1����?��
A����&}}��q�=��<w/�vso���'l�KV/�dN�T��4_2�1�4�B���n�w��y�%a���,M��gW����_��O�}���We����y4Zk[y���6@t
�D '���#8m��5�4]�p=��1ŵc��&NA\!��S:pi/���m^2fN$�#�w�<{XI�{�`���A��{Mj�2hƘ��_�b���:���]�&���2�����T�zů.6k3{`u=F�\E$�C\KйR$��`��F��J��.�Z*谪Q.'��?�S�(�6�9)\=�P���T���A��E��0ݟZ6L�]~��˯v���m�6�eF~[����	����!��O��s����V��s_�t�x령���\M�7���?��=w���EC����~$��1Mq)�p�?� ��៿�)RXϋ{��~�(9���k�h���ٕ���C�	�rߩ��'����zrN���>S)��~�_34�*5�[5�����4m�q��!� �N!&�[��u3�R9He�lVz�pV�ޱ�V@J4��L@`/�p���hHd&[���H��f�1�x���(�/��U����ΤT��C	2k.���f�/�7�6vX8ॷ�ң%s�MT
�]��mqѦ(�g�q��_QU\��I���챲��q�������{�j�P��
ț���o� t�?�sS&��W��-����@Hw��\�/��!	�5`"h\y	�3�{0-w�d
�@h�޴���TUa8A.��o1��v��&6�D����Y=�(0�EB�H��6�Z	|D�O��;�}�$p�ɗ�Ń�J�����X�v�f�"���� X�M6U�y�di.b���x�J�%��M5VCŲb�>�pӍs D���pD.�S_������ou�W7/O��
�`���6�I�>�#�	������i�*������t1[�Ǚ��V�S+ 3���:��5�9�辀���X7f������G�6����zP<��������5�)�Ɩ��L%\H�D`���eT�hAf�7Ȓ2��{���F��H��R�a�/�(Q5�ǳ[��=�P���3�$�jȥ��s==T/�WBc�gKϓ=��uA�Tj@���e%30v������Vr�f��#^�h&�R	bs�%W@CZ�b:�k�m�i�p�5C6��k�IG3���M�e�� �^�RC�1+`_7��hBs��R�r���<@f(��X����ڿ��S�Pn�����O���?��6K�;�Cu���`��*��.�Gpƭ���U�Eg{��^��G���"5�u��u���M��T�9���
�#r��8��\�g�v����ߤ�(]�o?�h�?��, D	��S�����)�����&K9�Yo�yU0������~(����_�Y�"�j�G�o��HGGMCO� �p��Wa �Ą����?KY�O`@:��S ��6�V9H;�%V��!]�ܐ�!4�B���t2]	JN�N`�xS��B�v�1+�oi8��e󕋹}�Os��*e��_vbeSI��;n�w�J,��������e424���"�W��9�G�[pT���qf���"_̀f������[����ച�*z�Ȓ����T2���!��-���i�� �V~@�y$
W�1�/�PO	��b
��V��M��B�r�[��L�c�%�}Ƥ�Q��v���5k2��u��	&u��sE�af,�ެ<A]��'��ga8��K"j�ek�K���DX��Y���b�	�/�gy<�)�Ծ����g��-�z�x>���̭�8�� )��ıEj���a���2��s/0���Qd���*�)�r�!}Xǣ�y�d�9���![�&{ж۞����ka@�.�~�ɗ���ֲ���갎Y��d�adR����<z�GXR00�HAL������� ��2������a�wN^v�d$_�:����|��d0i_�h��ӈ��o������Z���l�$�<�*�'k1�
��8���N�w��NzY�x< ��]R���۱?_�����J�Bα��׎��_72���F9�ۊ������:G�!�\GC��A�ͺ,�y��kwm���!@Ã�O�Z�FJ�:�C�0候�[����=*��mR���,��E�L����3ƵD�KE��>T��F_�6peO�<��k��w�h �ucU8$��pѭ�ֆ��}�)�v_'�gqʱ������v�(J�o�p�t�j��.�3`��uk���X1�|B�g֫�_BOn��	aa��Fh~�ش���+�Z��¡C��9kV����\�4N��Ef����j�C�9�<#���'U�y���C&�E�s]�h=>��_�4�<����3���e�?�V�6�y%���B�Y�h]���]�eW�S��w�G3_S�Z��6������J)y9����HLd�>_�&^RJ���t��:zx�#���xƱ3��^�?���v�Q����x�x��$�7l�>�"HQ8G ��4�gd����a�I>��0M�_f����1�F�VJ��(W�O�<{IC=�h>��H�v��qY,��nׂ�,�ԡ1͊��<n��po�T���xj�4Ŋ�סDaK3�
7���0$g��4w#��od:�{�X'�q(���W��Аɡ�����ᘀ���Z�IC׉P�bk�t
�GZb��v�2kZF4$$�渂�[��
f?z�4��oO=�4$gޘ��-�m��KYY�@I��u�5��*�ť�Z$�0t-��m��`0T�{cZ�e]����v�����B��}�wUQZ)W��F8LD�n�^|�[Q��$�S�Mrf$��I�m��́����a�ސPS�@�����LYQ�F��)��ҕ��N6SӸ*p��8�����Ovc%�~�a�Q� |��a�o�N|�%r�anհ��F�cf�X*1�϶ͥ�H��;�5� 5}1?�/[�V2�%��Y��}ئ�Ly!�S�!��zS�`��M��Cm�yis�{`3�]�{����R�e�S!Qȏ�����0̂�{|o%b�s`�b�e#�V�^�;K�$G]cO%1�cv�J�����x8#y�d��e���rB���@	������ r�ۼ����
=�Dw�Et��ǎ��Zꞏ�fݬ�)� ��]��Ŭ��L�^���{�"���������g�'�v����"As� �NH�
�v"���D�"8ZԺ,�4����v��s�_X��,�fY��G�r|y���k��H�Q���)y�*љv�=?�ɨ9�G�<)!�VT>	�g[��-{���橩VW�)E�Th�bn%{�oY,A�|L�,(A�q,��c��GVX�'�Q�\����:���S�#�k/[�Ď�X��k����� �Y\��t�B�[y��_����Zh���^Um�x�I��Hsy��c(���t�LB��%ä8��`����8Sh�֭0A�[�1���v`��"��:��ٙ�a���TA�,�c�/˾6_�P��Q��-ټ!_Ml���:{2J��5��7�aC��b���?��Qc(��+�ˡ������<S-�ͿG�5�׊��bV��A���ic�(�)�a9S��,��*@j��x���ΰ�*-B`�(v��
$���5ET,�q����O��A/H!=	��� ��_����Bd�����'&` 1f������v$M>�А�~&}V�Wͺ��`�x�4lZuQB���d*���3�R�{�J�D�)/�������绻�˧�ޙ|xLh
pr��<$�����,w�׎�D<���`f��/4����?�j��H�(IN����f���~�vzEe(��1�6�Pb���_~ҋÇ��1)Czn��-Y���ƥ?����4�j��,����Z �s}d |�.}Ŏ���wS�k��E���O�8�
Yǖ?2cͳM��׮v�N���Ҫ�f)�e)�=F�d{�6ͥm���{Y 7�\���^�>���������o��j�1d!���W�N.��.jA��6��\��S�q�-�2&���o$>���<7�F�|�I�@Zچ1�������.�v�rr�9��l�:�_��6B~A��>}�q�)<}z]h�y���4�(H�A��4.;^L����z�B�B�m�� +y[޴���\�7������-4�Ctd�F���2S���嵬�5!�uϵ]jPT��s����bZG��+19��O�f=3[zs��[��A����!h2��f� _ے�� . �h�4�-q�����c�f����_C��;[�KO�E�H��|�=�?��[��?Y�*�T��&;���E��?�Q��]cu!YIς���6��	u�pR�#ع�z#g�o��U���|��r�B;{�u���,�"�-�n�pGr�T��>�"a��p��!�F�&�A5��}��g����N�o p��2�\�8/A;�!-v�4f3J��P� ��px��R%�h`U�h�X�.no�����C:AЪe�ۘ�D���{�xF64�]���'��-)R��x�Ls�6��v�=2{jt6�%hħ�NUfK\���I�{:N��gA�_p@_*������0�O��هi��j�����W�Fm�''�5$G= �E�Sc�{u��"�����<V��zJ���&��D�B[�8Ѥc�f� �PWdw�H/ؾ1 �Ś_%�9���RJo�pV"63�	*��a���,t%��(nW�/QE�o�h��,�ȑ��:��(���ɩC��m��uo�b�
2�2��X�>���&��o��]�G�.�n� ��LN��	C���H(�oFм>�g���5-���g����~z���1��Ò�'�i	'���[R<RCi����@6�rk7�P��⩘n4&\_�S�[�`��K�PRH!I]�#��"+��#���-�||l�H3���r��K4KXZ�d�*;6/�<L$�
{w�=h�X;R���"��+]�v!Z��Y�.S=�Ɵ���ad�Gx}�`�&*jGΪ_�u!����%�ֳr�L��
��ֶ��ab��#n2k6�v��ڲ*�sLd���~m�c�B������H�.Ƹ�GPl�&���'��t.)�k������C����NxB��l]!B��=&��e���b�*|UA(�ÖNAf�j����8�Kt�J�މfc��lA[�p�v����G�
g��M1�Z�wXh����Ê��v��2M�X��߽ڤ�:� 6
��%nSO��PJגT؍i#%T7^�R�1oS�+�EH� ����Zdi�u�s����-�5�&fS*�&]�����͒��)��,���|�<�ѐ�gM؍-�9h�����s��j���i�u�óD���Zz2��ڰ��Z;1�
[d� �)��%Շ�[憜s7�Zk\O��#p�㨷=yf��!x�6D��e��T�=��