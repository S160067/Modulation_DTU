��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���,���`�Q �����6�͍	),�6�md|_��n�x�"u������K �5owJh�E��qڑI9����%,%UEwf�x����;.�9��p3��,/�֤����"��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv ��i��X��s�-�Q?F�`Y�������� I֏�׋������H[��9����ۍ: ؕ��6ж���Q��" ��y&���Y	6_���.���M�ݟ����k����
۷j	���`a�s�Yot1H���\2\:UƉR��S9w&��� E��s2�
Ly4�oW6VK�����L��2�$}�������H��N0�!/���%I!���G��Z�N�8���Dr�:$�B}R��z�bh��_`'������V��8R5Wz���ma��=l�I���@��k� }�!��P��*��)��ĹQ�F.3���cɛWR�*jN�6m�Y�ҟ�ݗ٬?�`����:��_�!�.�� p-F�d2�C�
� �i@�)�$�;���$li�Rҋ�U6��i�,J��`pR�@���@��\���y���r>�[Qc?�L�ez&��� �������أ��(*|�z�pƫ��_q�ST�F�{��[�c��Xu$I�KKu1C�D���J�4�0��I+|9�~E��~�V�y�\�������-e-��0hڗsB�jE���}���U˔^����I�AYugJ$���c���
����@j}9��!� ���_$���M�A��U�O�ݪ��lU���\�3Q`<�!�L����G/誩L���Z��ƴJ���a��!�I�sTm��b�����H!���$�*����%�f}���x�]a�w�㛚�M��!
dk����9y���i���c`z��$�] �nS)=X?�o�IJRC����8�(�\�r2+�H��|��̱��g�B���r�����K#Hv�y���3��{^�o�py�aB�DpMZļEWbg�!R�{*�!��|���N_�����s��Àw9������E_;�>lU���a�����|��s��(q�Co������ˎ{B9��Ķ 7�pZ�[��O�d�q��Z)�+��z�����E��V��>؋RD ���򌯂�:=d!��0TP�;��!�-|*Y,O�-�8Qx��Z��K�_W�7��J_�u�<���u,��[�Gf����P��|���7$X
`!��r�B¼�R ��J�]B�^l�k�R�WQ����ߨ$��e{���Ƈ.NHw-v������a���)05c3&>^L��_O���:ڎ�[�i��s�����E�µ\�'8aJ��Ҡ��՞η4�5xbHhG&L�{�k	��P��O�ޑ(����pӽ�/��D*�����E�\���Hk-V�ZY95�3�;�	�ڬ�[s:��w�����p���@�CQߖ�b��R��u2����r��7��!q�����ДȜ���\�lx�6�������
vW1�&|R�m,܆���>P=�dc1ѱ�Emk�@f���`O�M ��	˚ۢ��b�Z��.cޤ�{���+GR)I����"c���G���aN��&N�K�9�Հ���I��7�V|t2	k?��Sf�0ӹtFGN�&	a*Qcu2����[TMNz�d�B�F� ��F�2��/`-�n�~R��^����$?������ˑSvǃ��^�v`
Z/�@�n���ا�֧��L�RuC@� �r򝈬��M"��m��q�x�D�H�$ܭ�����n�"N#�AV�g �s�I��MM�0A˩L�z�G7f\�7�fĖH${�&����sK	Tg��`7-nó��!-/h"��tC�]���s���&����Q�?�$�A�i_A*���!�#\�	��q>p}⸫���{�,�;�,+h�x�C�D�x暋��E�Y���䏮�?��fT	��	�����̅n�/H���w��9%[z��rQ��و��67�����,�S�)�n���+�d=���ah�����&BV+�T��u�A1l����o�K��f��E�/����2Ϲn��D�gA��ꁦ~�@�UO-��o�;L��8m�cn�☂2tl�����N�XҲ����O��b_�ɇ�2�-O�+��l�����T	�26�E&(�`���% ����O�7j�ɠk�Y���;�#�U�����
̦Y_��!�G'�J��2ҟ�~�Lto�Mv<
��o��N��6��#Kն)��F�#CK^eӎ��D�D3��D��`�hY��u����?�� 2�D����e�?��>�Ǻ��ԟ*#�Gh�T�/V/:�tv�J`U'���j]�MwU��q֯B�9ב���!� JʅC�&`�u�$�b|r���3��FuQ`�����32�d ;��b�Bפ�5�١#9☥��A� �:�{$�!.�$���:-F"����cIR���������&0�Čp5��K)D5ѣƨ���Q��|�FJ$D(s/xt_$1�<�$��!�w\/8�� �i�XR��sH3��x=_c.��+�gT�'<y�Qҷ����)'�/1��6���[�:s|/�7M[�Z��3Kr�b�i\�>~<��&3�����Ï��9q����Z>1�D��9�O)����Ɓ@sW)���w&�*�����j��. �0h���=���8�Bu
����;�^g��A6V	֊�鯨�L�2��`>Q��}�x�� ��f����V��<}@{�;��U�k���_(Һ �����L�SG^�/x�-r��v�!�~���p�����f]��k{#��K#�ZHrh��F��	�O�=6����p���Q��M6�[�������.�bE��5S��1n�l2~�#h���Gܷ���NjN�~�VĤW���%�B-�Q��RΛ�� c�	��W�
��g�tVivU� �6�K"ޞ^[�����.��|�<C��.�i�ß����MTt6�@�Тe����h9�25�.���K����b!�
�tdM���l�M�&EÎ�4� hR��')mj�+4 bG�j���+(��&
5�%i���ma����e�:�gs*�>HX�`)�k؞��$�2���$C�2v�G�`b�gx�k�O�^J�{�
���	�w�Xr��x (����l�n���ӊ��%5��>�����nN��C��O˞|�=�ao��s�K`RY��yUk��\z<*��9|�	�#7��'�$�Ka�#�VHB0C.��t�/�����,�m��88���U4����:5NDyn�/F������/02e�g�a� J!�@4Eg��'�p���"_'��������o�eP�(6�:7�L����s�	����E�*�->�a�L�)�Nc5j�����H�b��J?w����鑎@DZRR�c���Hy�b�"P ���p)���ߊ���XvgGF _?^.Φ�;���~F�	m���`x����M��f����-�Ί ���_�q&4t1��|�Z���h��F����	ƙa,\"Rf(POI��D.uoL_
����œ��P1�C/Jց}��]��A ����ff�fۋO1T?}���Y�(�R"����#���"�w��4,��=���Z.��Y�;��:S_	1;��hO-G˝kt��u����dGQ�$u��`��@�X��T��>fh���j\X�`1⊉��BbX
K��Υf@RoE8��9q�@tg��������p-Ia�Z]`�%���U��x`>�դ&VxP�7���Հ�Bt?�i��� �g���0d]{��z7�7�FK1�5_wdb 8�?�~.g?z�S$�ǜ�s��2_��岜(}c���6���h&�LR�1�|bK��G<��ߥ!�o�=��c���z��Lm�qZTT���Y�U�=q��%����}RFAd&Nw+�;r�%���:��m�j����V�ƶS�ٙ�����*�n��R���-��[qJ�}a��ĝ͏)�JZ�Vq������B��TX^^��,��A��mF��c}�
7qcSj9l!�GNu.ӏ~[���<����9��e���%�y�b��m E!�g�^�|�������y��A����V�2�As���*;��/��l�r����qob�	x�
)[�!k�t�A��!����J:wД!i��.���"�+���	ᬵ���M�d���t(��0��Tα�������#�JO4|�-��I�쩱 >{طi3e�q���Dz��Y�1�|D��D)�2������faWe�%�l~�Vf�8R�7z����u���ID/r��}����tM����f����^;O��3 +�GNξt���L���US�x܄��ϸ�K�A|�v���y8Mb"�KŠ�P���`аVjjW�I���LD��ղ��&��jղF Z����PgN�jY.v�CV���k.�W@�l�� ����>�d�J��`����T��0�Q3~�V�r�:�14ц�G(ֆ��R��N�~�K�2��몒�ݺ�V�˪��'v���ap~=�X����b�yJ���<�9����F6�%"�#��֍�����?��� x�3��b�G�/�����Qqԉ�z���'\��@�@��$�}����[(/�9�r������_�O�����#��4���@��PH���^����ɲB�ԉo4�e���$^��N&34+� T��9���Dpe�5y�p�/:(����`F���(_�*��+���E��1��T�E�@o
po9�>#�� ěK߅������,�¨e�"�q�wu4� �Ze�1CO�(�{=�pY>�E7r��sO,�_�
e���S;vFo\ճ���@�
�1Z�+=�Z��c7����r#c�_-��wƊ�2���DH;��"�XZ�����ߜ�P:W�H����[=�I��B�,�p>����c�@��K-��KL�f�%�m��pse��v�� j0��!&kз�}
�^���oo�͞����ه���Ǘg�pY��C�;̻�� 0���
c�c���[�����#*X焢ϝ��������%N��i
U� sB��%0����2��?�C���J�i��O{vf�x�zQ�(žu�n&d��(H,�(T����:����'j5�R���ra)���_�M�̞�bszMմ�U�m�6�.�e@Ks��F�<~�������{��-�ߟJ��K��44�^��?�X$J &�"�"C���@*鼧b�� �+��rY��Nf;X�C��u�t�ߩt00��*ba/�~�(M60S��#oE+����N��x���p"���)�
=�s��;���vY�~��91[(^j��J��j�l"��d�]�;��6�6/�~KI�qn��K?�\\R�0��^ɒs�<g7k&���΍�偻�Q�5�~�2� �DT<�B���q8�|�Ag$#���7f��<%R����񓘨sJ�ǀ��Gf�M�D>��=J��1Ҝ�,�l�]?��/�<n�t�UQj�8�e�P,��̌�h)�*H�ռ�8,��yN`U�|���Qr#�x�GYP��4�� ���/GV|a��k�U��=��m���;�m����c��21�����Jv���B9�-4V4{"v����̏~uف�O�!ͮ�g�C�q�����j�Q}FP<�S�9<"w����<3���.��r�u7,�1ˏ�v~������	�6Sn���D������ܨ��K��ȿ,:�N%
F� I����QF�:�} q����Ͻ7����DC�g�.p����>��C��{?[l�];�x�Ч6��c�1o������X�vV�e����C��l�R�R�_�U�%墕VK���0���GT,��,�S<2����7#լ=Z�?�(I_w���F�ff%m�(��?����G��0Wp�i��O}��YY->z["W���_���x~K(C35;ג*q��>�J�ߕ׀XԶp�k>�PVMI���LJGa__��q$� y����UH�۱1��Ք^��b��e� ��1PM��Y���V7�M�zR�QW�Ϛ3���ˤ�$�`%�V���z��V�d[Ms����Ģ�($��GD&���J�o��n�{#���bZ�a��Tmc:�K��b3]�=y٪ϝ�5�o���ޑ*C�J��M����U��Y[�K�u#�����QYV������k6G�M�og��2��;��>���XX�R��u���L�4wt�u��ZVC��xX)��[p���y�������zQF��rng�����E�O�o�Ԉ�fq�ӕT�%�[�NH����Ht/�g���8���� ����,��/��`��hfw��f�JЪ8Mz��t7���[r�f�{hQ�4�^��g�c���
�����-��5��x��Q�$��*�r����a�	����e&%D\�8�jM��z���zo?}eޤW�E	�*�^x��N8�ٔ��u_*wR�#X0���/D��@I#�Ͼ^��������]C�G�ڜ��R������Qr�N&�����:����uV��,e�r�i��
�����YYw��b��ԋ�*�e�+U��|�AP�Qϩ�p�R��v?̻d埕���6�&��<Q�HÍ4cV���Ǧg�3�'��!t��-D���Lnt�ڷ����QǕ-.�����lO�����J����" ��r篯�np	ReU��Q���wy�	!�+�T���w	� 0��� ��9����R�)Np�-�gHis��Ce�%���P��A���n���bԍ��"jr��j�\?I����?b.x(��Bh�᧳ҕ �q�����F�;���!ķ4���<+o��k�A���#���d�<kj�&;d	}��������P��2k���[S��z�	�ka��?P�uVZ��j�9�.�cp���1^��`�/b�Qw^��U����`�N��*��b��0�� �5�q>E�1�)�G�?��|���1�i�6����;4�Dσ+����\�|L!:�0�A�K
��៶�4X8JC����g��c�{&�(�&�L��7�g0���p8&Уz����O?��H�B�ُ D��m�-�p	�O�8���~}FX|�V
��C:V*#v5�M���J)O=��z,Zrɚ�M��97�ޟq�V�<���ё�#�Q�]�)��ߺ)p2DR�lnY��9L���fdY;�3ȁ$���lo?��P���YXWf1�a`���x���`Ĉ��;�G��f�t��)��N��e==y)<S�Π��m��HM9��&8�B��.Iҏ<WR!\�7���^E�r����K��z���̲���&�i��(�+\߼�Zv�հeU����,�����5��K��o2��Z������x%����ؐ,/Y#:01�l"��ƖX����/B~RҴR�Ki7�{9��&����k�x��u�IfsN^b�%��Z|CsrU���<)��\�Da�x�����	(}�Yp8�ӛ�Us�|W��9����ӴN�%�W�3$T��G��Ҽ�]�U���z\��Bp�D,�f��N/��=&!ͧJ�Wf�Kiq�q6-��a�1>��X_��nw�O��e�c��]/���$� H%'�(>/5�t���ג�|]�gY�}q�G���IМT�R["�B��Y���ht`U8]�uIfu�?��9�'�ʶ����	�J�H0�ن�̷Y�k��iP��{x
��!�ϝ(�>�HDZ�<I�SA?�h!�KC��Ιk���@*��)	��!��j��P���x�f{�pW��x�dk�ـ��i'�WWj��[ܛj岩'i,�e�9DoA�WJ�8��\f��W���
�����u��Ō�S����1?d�����U� t�.�qՍ�n��܋'�^�k��'�Ra�-�NGw��o�ͱ��4M�H'P0�4�
�xfS�9�P�9r%U7T�#���$�H���_w,�N�Y���י�
:w ۣiҪN��ȑ(@��i�I�ٚ��6��o:��:�\A0n����
�v(`�?�Z����#������b��sMm�3��u3�*�W�O>_)��L��}S���3Bt�}j��pgA'�HL{DC�N�1̻7��ܭG������o��,�$a��-X�ܓ"≫8%�@�c�i���љ��y�2刽�!T�n(�#9��/�|Sl�C+6&�\���	���Si܌�]~�suϮ�uwI�����T-�}hT<I���-��)�L�Ι��H{59Ŕ���p�*�,i/�D���*>g��
r����x��Kݾ��%g�C�D�!�U"�3Y�7�`��B�sA�R�>#��d����b3KP�gPLWfV� ��5�L�ڸEJ�1Gc>�՘�����[������/��	��m�����Ðg�~����N_����zH�z"��6[r@Gg1�4~(���K���U[@��}�{sS��Vd������=�^��:���*P�����bKYSmߣ�8Ԙ���<�	2-|�|�`��x�K�g��e=�g�\n�A�+�r�U6�=Fm�W�;%��\�1���|P�[q��@m8�����y�8�����5<�^TX�/��7�pOIQ+�Ba��[�@��=h�}G��p�w�=�tx)�i��g{[���5m�p��y\������%�N�HoI��ӟ�d$��q_�.p�F=po��Y�B�s�n��G�P2-?R��q�@i;�.g7^�4yi}��v)�/��j2#"�rU�t3���(��X.e�W����S&u������d?I���:��V0�R��-�Ǖ�Ѽ�pk�|���x�#I^kޮ&���	57}�2��Ao����������b��81���pL��w�!Wx�_��VdI%��i�o�Li�@��������^;�,l*|f���y��x6�[�n���� �p�J?��p�nMe����?Sp�m�����������D�&�l�(?��'ra�Y�;̎�����ȍ��n��Ieʫ�	��%^�8����VY2A��t�(�X���v�,y��U���ZXֈ�Β���{pZ��_)�x�V6R(_*O���=��;���G��I�|�%�v=&�� >��&��.}B����d�2WO}��R�kdˏ� (3�F��$�h�D��=}w�+!����5��3"u��|�t�"�yTYM|���ćta�8��u�i���Eے����u]�QlW4�M}�U~[K���������u��˳���kh����ũ{<��L���L�P��x�QX<QN�`��� �<��7�T��jk 6��!��/�.��-�'�,����QC�s�`��Mi^ƿ���tc�*���B�߭�tHC��x�a���ѐ#P<���.ƈ̬8/-8��?e�a58r�"���Ք�|�m��y��7��ilU*��7;��ٺ73�xa7r�[��V���Οɒa��7�l<t Uk�'jT_W���E�.�d��t!��5����������Y��8��YbO��
��C�#��f^�{�����bE=pUr��6?,g(`�UG��\~�!@�y5��VP�.�Zk��E;_������硏���B�$l��!�yn7i�a-B��m�E��H������)�(C�B�G]�l�����ģ~X|$L�5@D�qg�?=�6�ķ� ����Zخ>B]���L5��f�y����:{���/UnF��Μyƾ��+zAֻ_e�����:>'_Q��m`�r�!L�z�[F�lr5��g6;λ�2�1/1	J�L�_uG\2G�|Jn�G��������|ᆲ��]��U���Hx������/�R_$v- ��4����j��H�/����b�F�3Q���wmy�G�K�XGĒ���tl���R��r�vh�?���ڀ�:�[���ԍe'�sw,x����S;��@Hc}n) �4J��h �{=z9÷l��8�!���,jt�PH�X.~x��}�
x����M��F��ĭ`)��M赳2ǈ`��8�ٻ_�ذ}�D@�F�G�-!�; ��)�ǎ�0�q 	�t�u��w^�S��q�y[蔾��lq]����Gry�� �U���h���m�m+�l�5��]���59.vE�+(�^$��*_lS�kŦ���(BK���J����y@��>�������Ы��Z�o��m39KK�x)`��aW���Gpg�*ٔz��FBD������qCM�G uio+�a;��A���G���X����zT:D&ԃFg+i'�0�ʡ�[�X6.h!7��/���4�� �0ܟ����.�y+�q�n�j�D�}Aa4�����Y�W�[��7�B/<YI.�C�
*!�k9�;��D(n�Ɍ�S�o��W���#k��XΉ�|^�Koz:�c$.B��:n��&�^h�9���Y8�O£����)�n�0s����4&��X$�-�0���Xt �#f6aU���Y`ݖ���ƇH�S�>֬a�'��3���� W�J���?,O�_1�L�}s'2Sh��1��+��yۢ�0���� �e�z�]�&���F�	���M>@X����;�w���>��'������iCx��P(����_�l+ꚼr��}�'}�ͤN�ӷ��:b�LfL�J\��8�
Got���7�v߰*��7�JӀ��b��h��W��V�����V˄�I����\M�j�����{��S��[��M1�����gL)	���">%	�
��q���%7/˻
�t`d���k��8�L�I�)�V��7C�d��sȳ��j4���7�Y.ׅ��ي���q,����e�G�|��Z*�_|F�{?�J�ɱ1���"����Wo�y�5K�E�f�����o4+�̑��j;��m�w��.��C�h����[��S����pJs�N�δ�v(Ã�d4+�|�p�/:ۄc��g���{�࿇����:��J!I|r�������ۋ��,""�n2ht�J��5��-7��O`y����9-��@'�L����o��)A}�Ө�)vS�� Qǩ;[�w1����ڂi�r���*����ۂ|���L�U9�����,`.��5ز�0�ìU���x���D Og��������q�͗���Y����>��E����&��N�j��ŧq�ŕT��VO
{�����]2�e�T�K͝�_Dm�K����R�=kŴ������гz�{�Iγ���  2�c417�`D�xU�K���`4:��$>�� SR��(�W�yAB&��;LF��Z���}���9�&v��]<m�Wó]h�D#W�1���!`Pb�k�*���ʛ�1D79�|���R�ᮀUQc��G.���|�O��C���k�u5�l����w�*srr��Q��IEae��D�w*>_F>s�2��h�o���ĬV�CT�|�D���>K�L�u-�e��O[g�Kf ���Z�+?m��]LU���T�gR{�Y;�+�nݺ��`��&��z�?ӷM.��z��́��і!��_�n��G,�Y�^���ԈE�'=s���6��Q|*M��c���*�A�fH۩MM��?�{sg+��o�9ow�W�_��a�â��hWv]ǅ���xR�H'h��� ÎG�f�d
���o�~�
���G%t�4���7�/�2��=cY�S�3��D���51.��U��Xͧ>�6-�p�3ַ�+W���H��a��f]?����B�ި�1���B��zݮ�M�A�`�d`;^�y�;
>�/��V��!|8�P�R���&��r���z[�*����	��
�]Vp���5�O~X��r����г�)��]�|ws@���ƀa�U�,�&�vq���=��"Ŝ�!�(�f~���cn"ԃw8�]�?3�Io����`���p���^|��p%�oK�#�cJ����h́V����{,Y<���ʿ�Y!4���A�����6�� V^Ʉfd��Y�T�̭�����T�T�)�p�\}��m��}�Y(p���oq|%	_)�D�״ ʧ͘��� 	��H������-�ݖz+'8[��v�CRQ!�('�J�o���5��#�a�B�Q{%�?@�rz3'�>�T�A����ᬲ�b��5WR3WQ��:��4�*�⾫���{���y������Y�� ��Ⱥ�Uo��."��6^�V~-FI�U� 0&I�`���*�B�<�T}���Uא'#���zX�w�([#~�p?��(_��]\��1{�[�z�j����5�֣�8~�-djaA�]tqb�����(8h�i�H�5Ph=]�{1��}��� EI�ّ��Q�zS;*��hu(�]������b�'Ṕɼ�q�H�X�1�'��ƕ�$�3�&Fܘ���y]���a�,Pg�]�����3�󬰷7W#+�U��4v��=��fȽ�~�	6���P�Xٻg�s�qT������q��z��}9��i<N�g5�r@��=�3�R�و}<�	0��q�gj�vu����qL��`���O@\R�ic�@�DM�/�K�4�M�y�H���������,\�5 4����#m寧X�y��d
�l��^<HQ�r��ˢd%���,�.
IT��ɱ!f6~���Pcѝ��ea�txJ�#���X�y˖��k}�#؟`�����/�K*�W��8�n�la&'�9������!%��9�5�rt2]��-���W|�A�
�M�y���d'�o��Dek�栱g~���#A�wE0~92 �y�~�+s�����j�W#$�2�>m,i����\R�������r�%�QS[��L�h���8|�A�{ܛ�(Z���Q���5@�]�,UOH^�$�	��"Ϭ��44������4�3��v���� >��%oɿ�h����許�f�5|i����L@���j�����ҧ�����Pr�"_>O_��I��`�0�5s�`�g�˶0�{5m���H<�[o3�O�
k��E��O�79j>`�Q�ލ7@W�{.8"���}���S W�X.��v��ʊ��=�0ep��f��&6��r��!�؃ʮᰌ����rQ�q.+:]�Xyt��lM�cV�>$�D��h��ßNj�h�,����qG�GX�6�0��8 ���5_�vݐђ:������}!-�:�r�?Q�(y���
/�;pą��׫�5m�3��;K=�"Rݪ�����٭�.pQ��Z��ï#_�ˍ/����aA�LQ2�k����Tr�.'W.1�r������cK�Y!?����7BT���&F�����R}��k��_xT.��Q�)��?(�DSU)A��H����}U�о�F;�;�H����h�VQ�niHJ2��Q��C��LY$|rj�-�}�ʼH�'��<a���/�0cK�6'���dp��:�-���L"}�e6��_�TA������]����R6�����*�>��5�����p����`m.�����=Og�O��1U=e	_�jCT����6VKM���#��Hn�#����"��/՞*p|0�v��L�S�˞?�v�:�����n$:���x���ؼ�6��7[/ԿٵԹג68�:`���˩'v��:_�1q�<�r�G����RҫX�|��SqIZk�V���`���(�u)VP���Z|_�e7z:Kҽۋ�g	�ŊK�0��k+�Ov�bs��V�>jv?�^5k!y���W����R�_B����;h�{(�diX1�n�ȥ�n7$��wqVx��E��7k�;������A(�FϦJΞ9p���:�@���p�9��B.��ŃHLv���)]��kV2�yҾ˔᲻Kw"�Yz�4OI�P��{W�A�>"�7�!�D�(�{'Y������ZV3�b�T0]�ޑl��)�S�Zрu8}�c�:>4>6���"��Y-�^k�[z����dH�%������x���;0�������^u���{��:׶��.�(�S�At(���yJ�E��'�Ӯ8���ÃÇɻ夵�W���ϠK�����[
���Q�?�TF,C~��>��~� �t�1����b�����48�}�h�:T�v+Vj�W�A�f���+�	�ͬoV5E��S�F�{ō�.�5��L9�}��kC@U���1����� �*�D�:�5�Z�`�L�U�_mb���$m�'
��z�<)�>��S���[�G�@hj-Mkjٛ�h����d�������+1�<����UʟF1���dv}�6M��p��Fg8MzM<Ң��>��������[�h�LUx�pǸ�V�K�ZL���<rwl�����$QS�0�	����cI,��������M U�ܞ=��t��2c�|ѿ�n2�2�+�Ś���T{�N}��c�U+����yn�����N��a6�/	������1�,���G+�4z�p�Sj�'3!���sryjMw��c΃���"�V�`��y�_�9^���o7S�m�w�p�Y1yG��X�ִ0���-\���8��-yD�x4�����P#3���)b���hߐl�8};��pF,�ucJK�%UR<���3��av��7g��r��^���12!�Ć�t:3��2o����H��E�킙BNP�����#$VK[�:{��6tX�J��BN��3jZ!fL���.r�կ�d%ޜ���I݂��@9��T|�F����[;#F�}�!q��;��3�	�~:���ĥ��ꐪ���lb��@hW7�z�i�z���
2��]��Z�,	�ۯ�Z���$i6Kv	���Vą^%�$f�(���3�>�i꽪π �c��)V�<�K��M�z���چ����6^��"�SԚ`lېXV6�y�}��d�� 5G!]f�A=\�KW*�8'f�􃻠�I�@�+��W�������m/Ⱦ�j�O,i�v}1�G�c����¹/0����W]���ג�����Eh����8{����Zͩ���̩�a<��%t�tfI�[�@�B��	68<�R"�Ӥ�4R���^hD�p[]8�>�H��mS%��sw�plG�彿�fx�p6�e��j=�$^����9��⚑�x��7=jV��8�y:���ą���~��o�yw�\���#�u-;w�ey��ő���)��S���b۽`p�5?�Z�>c爍Ա�H�Z��s���w@s�g۝����R�'?�ц�٥T��u�c0����<���ƾx�La`�
Q0�k����{�� $^�Ǖ���D=��;�ׁg�5~�<`qWT�T�}=p���7	tg�\y2 ���x�2��T�O���}ޢQ�6�`T{�B#k_�
��}/���!ıK鯗�*84�l��rHq`+�w��<Tڇ�*
?b��1E��,�]:��Q�MyX � lI�����\f�܋x'*\�X��*�o��� ��j�A!-�V�#���2���>��CX��>��&�i�wK�='"P���*�2�]߆���;R4���%���y���ac/�̭�����y�0y̒#��۷6��R�v�>	9��n.�C�KY�0�z��SiZL#��Ӹ�eﶔK��'aH�ZX��Ȉi*-ACY�T	-ޘhQ��K��N�i�ҿX�#{�g�uif=؍�nR�`��n��XT&f{�LP����`��6���Q%!��0�,Z�k$��N�\��U0�seq�0�J��m�?���Y�8��G"l/��� ���׷؞F��wr� ��NƯ��@@Tg\_�F9�vjZ�I�k����6��At>�g�Aӳ,o��!Qȣt:ZCG��ciS����޸$?�+�fs�Gt	Eyr~�#��|�i9p{��$#���'�#��=�X&��;������{�!D�?
i4��G�g�0��Y�_���� V�pg�?L�=[*�)1y�.t792<�vwY0bl�R��n�N.�o�0�꒴#I�qsT.ϚLq�q��R��FWUm��٨�r�4�*�mV�8]�ZD��2�\duW;,�m{/B���\	^��|�@U����la.�9N���;���5�|��;#G}}(N�(��ے�bCWp���K���o�pt�"���vɦ�(�s���kC_���
Vb��#�yť!*���ow��Wa^�Mx��M���?D[�]��U�f�/r����i��G���in�:��ӗ��] �����5�.5��ENA"��X�{0����g�lpZwUA���a4g�"�>Tp���b�w���|� y`�>�](6�t�J������@�}F� �&�}�����|�V���+��ޒ�ୂN2�T�������d��<��)���(�}�/��.����&�"�GW�\�����F��/;Mi�V(낼<ļ7��� �#�o�����,��'�E��b�ce��' �J����K�8ܽ�:����p����;s�֚���sj���f�qw��Y��{�Jh=V�~�2��.�gm�z�jBR����������U�;�E'�����-k��~!��/�aB +	s��J��K���M\��,�sÙ{�:�j�/\#���u����"3/�TҰ��~�&9������Z�5��Y�Ka��O��=�R	�:�<�����b.�2�¾o�|S���^�έ&2GQ��t�@�sэ���Odn�ͮx�CҌ�<0zP��_��O�T���\+ؙ@��2��Sh�al^�_W��k�N�t[$M�mg�<h�M��#WC����^H�5w� k(f����MF���a]�RW�,9z!�]^�;���[.3�>�X�P1�?�C�S���r���sp7�d�qp���ן^��`�D����ȩK����u��bfy�'(�v�ojL�(>�ߴ��;t���y��Y0D'@�uKّh������I�C�q�yF�'�F^���~Q{[<�.Y����43��GL|#�P�Y���Oy�Ҳ�I��9�b��š�l䯗1"(�W�C�^Os���Xep��'����I�1̢w�>�)AX��ࢀL���g�N��; ��& *��y�!��hވ���@��9�c������2�粞�n9���Bލ�K{q�	�����td!jq��l�e��B++�߈���T�	��(N}7kѰ%����`�&������x���7��x��^!6:�_�V�oy�� �K��F� �^��|�ou�
[�]�E�b�X�~Gh�)H��I�qӀ��F<#}l��Bӵ��0�73>�� �rrK�P��ʵ]�Ğ��>��l����"�s��r�&1!��*��o� ���Ս��l|+�˭���P����	is+�V�^0�Zk�M�B��T�0��-=M'��Z?_�I�����֜�ӛ�gi�_I���_D�̢�p*�I3�F&?��"$�m����:b���e�?����Ij��]�h�ӥv��ϖ��DGB�{����lH(�^��5�R�.������z����ˈ��A>����t��w��֦$E�(����&��a��-$3�Ʃڽ<<�������.ꖼ���;��y/�β�����-�.Q1s�]�͵n�r��$�ҟݙ?�e��6̧}`�5a�N�U�Jy���Gd��P���09������M)�ʰ���5H�� � 9����p�uU���ӗg4���j\	�y
>T�7u��"��D��zh�� ��I�yjXM�w_����g�Z^c!#P�^��ݬH@Ct�j��{����g�a�X����%,�
��k��h���H�y��kg��.�nS����L�E��q�@՘�'�����	�^�rg�*��7�^L[?�<X6�0��4��E����[rt�#�v�q@Џ�A����$pg���h�X�N�C�h�F�BnCd�ܻgmKa��Ǹ���ە˕�K3�8҇�])q�N���Dt9yި0�Hk�9��@[�i�pτ�v8�*�����������	�ݓ`B�ÌE7��
���8�L�Rhe&ΐ����y��*\���v{̸�5*��
N��a��*��;'�H�:�̂~�)� �H�>V�@Z��{�6!��X�0�����-�u���:G�Nciv]�>&�?c�b�'i�4̳�03�91~���&J^���s4�Ψ��Z�� �Z�ihO��PWO,�W�Tߺ鮚]φ1�(�P�v��\�������h#M~��Pk�ym��?�,Y�Y��hb�Y�.������8Ľ*�K�'΁a��J�[�8�;u�Z^�+~*��$cݘ�@5�:sb�v8>��{Z�s�5Җ�pHlny�U�w��
���U/���\�;oY@U��|�����9W��!Ȫ�M�j�"T�\\QK����~��m,KV5
�
g������Ȕ��� *`���{�;�q��X���"W�*+:��@�[�cv�Y��͌Zj�:� �H��a�-�>�m4�o.�D,� l����f�d��5ǧT�`�&�4&_d���&1���p�8n&[4�3�)M��w��J���c"]��iJ���	'�H��X����?��\���
�\���i ����3I��سЗ�W�&f8�:����g�k[�U��ٱ>���q-�b�7G��)��n��'X�Ț�*�e�b��O��,ZDN���/�b���:'G�B�ț.���-i�p����Jţ��5��h��m�'��+�V��H,T��S�&��1����E<���߻6�^�͍7x�K|£� z@�o��+����{o:9ܪ~�o<�'�����H-,^L������גmu�~��%�ld�u�
�Lښ\��1ʝ*=��O�Q��>#� 	�����������r��?��e)s���o��0_�&�ֵ��q��u{r��� ���;Z�)=�y�vx�z�c�S�L�a�b���?%m�0^�E(=�����ܳ��StC� I��<���᥃ßqb*ìy�xPs|�g�K��n�stM��K?d����'.���O>Z�'͘�i"�ns�J���V�ǖ�œq�L����芌�z�E��
�O�?>* cso�2㒩��`՞�եp�U)����UX��=ژ�ZE��4�{�ׄ�$ٞY�+�R��##�O�<��V�����]�?��7�Ѻ���,w�F��)�c#5/T�>�F1��-�eBw���q�+01���s�&d+F��`+����E���o��{��+($@�tѨN�l�9�!L�َ.��B�'���A�H��[~)f����ˆo$�5���n!b�H�Qa!�6���}D�׊�P�q0���c�vITW9n�1E&�H��e1#�%I��8�Ίz�/hG6R�͋È��i�5��H;����U�#�5�U���VT.�b��c� Q�����i]����Y�!D�$*�i�*�(��[{���9��iG�����q�E�"5��«&_�$�u�5�s�5>�&��6����])޾��ƒ�!L[�T�us�	9����Q<PPKj�-s��<��{�i���n$aR��T��24�B_V�
,�j�D!9�&(�O-@�C�@���<ѫb#��B-sQ�W�5t�'9��ʒ��"� ��Fʏ��%b{����3�i�B�&S���_Pd����d#���3P�� ��~� ��2��/�W 	\�wǟ�}�v$��~w{l���Ar�ISt�WHj���as����]�}Q������uGN=z�]�׳T���YI�|�]_P��cK�b�Q%kJ�-�˽��޸��C�45(8�E]�t����4�ZF(�����K&��	*qO`�^f+4�kG�������9g<l��c�]�Ù�1s��Fv��	֎��à��gkB#�K��/�I�^1�y���`z�\(^M}Y8�I\�-��������un����<�-=�:
VVP��Z�������,�wpC�}�R�ߑ�\�[TDMG���9�+3��C^��ߩ%���M#�E2ס�r��]4����Q�y��|�Fq)���G�R�T/��������g��J��MY�7T�#!�ȗ�;��l�0 �S[6�:q+J%�Yؽ	��.
G=��ki60���veeᗔSy^t�$������ �-�H��f�X6.���@�PQ�^%�P�X��������3L������������I9�a������c̤;���LR��1E��̏���T���߄�D�՘=z��V�,����H&/����X��7Tvِ��q1SJ	��O�׆�_ \qp�g���2-��*��E��������%�	~]�X�t�I�=��M"��}9[U~Dj5P��@{��ݲ7ݑ
ţ�]�`��Xr9`=�sB���Gw5	�pT�&�q��mY��1�.If��H�����'�3��'�6Y�$�|�(rO���%����C�֠Ɨ��7�$rM��9���P�6V�z4S!�}>EqN�0���1� c�d0��w�Q��K|uӉ���U ��hu�u�c6 ���6��h��)>�ފ��x6lX��&�������C|�Z���<��Z���ܭ�
��$�%�"���'�0 9$�nrQ~�-�~z����P_1�H�*zouó�|�����QlQ�"ם�!-�S�'P$�T��m�e������[��P�;�)�4�Ѱ��R	hB&�,��c����A�Q7¶4�����n��w���X���������`M�:l�m�cp=��@2O��ϊ.�����*:w��Ɛ9�Z��/?H������o��NK���bS�(���8y���CI����AT�k79����D��}��"�2n�[hCsş#�u���y��R��5�[8LC�Ν�b-�}i�s��V̥�
{���E³�o�[_���H�ۆ�����%�5W?c;{D����63�D�/�L�e(����5.��l�឵�.��6��9��>���+����W��:F.?1�}@(,]�����=�B� GO���<X�R��l�űpG��^�!������l��M9���g_ bg�S����8��QtJ�&"�Dr�W{��U$�F84ϟK~X��m�P�<�����)�>�*�׶7�+Υ�[wX�(ņu�k=���!�� �ˡ�BF���"Z;�4���^��bt	�R!af�k��>�xFn�~��&�K'S���ݠ'���h�7F)�;�F��9�I�5�qD&��`�lܵC�Xf������'�ǣF󯹽:ɑ?`yC���̈�Wqm�3�1^������f���(�ͥ/-�:L�8��ҩ;�5H��H�u\�j�WZPxPe����djs��k���gߜ�2?��R�f��/-���sdCd�N�2�m1�$�s��nޗ����/|<h���yO�����_  ,P�{K�����Ycs�Ж�ۼa�}����WW�0��I$�I�V��K�2��ӵ��8��C�ww~<�΃"r�c��a�ɶxģ�Xђ�˾���x1�x�\9AM���G�"v�ޚ���a�ά��O��j!>�+|^S����c�@��kHئMc�="@�Wo!�܊��7dh�W�uy@Dշ�R�0��Twdy?�Ad���D��� �ĉ����}�܈X2s��p��ӂ�x��=Qc��l�/�Y�JL��W����ζH�i��z����eh�䟋�u�����E�z��u6��GR�A��U���3���3#�p6��L�E�W���
�~��L��:�x1a��يi�PX��^*��8�<�6]�!�?�d���H�Y�i����͓��d�n�#&>/�W�G�w$
�cm�p��3�M�	�S�F7���)W��#����*"˾�C��\P�FGu��-!��P��YF�C-}'��c-kf����~o�l�A�O�;K��*0t�_F�[�oY꾳�~�Ѧ/`;�<ub*+���j;�9.���0n��^"�n�@��~�����Q�]%f���ш�(T���=�PA�{�X`փ��MGL�W>�.�&����O�j�g�(�w����b����F������%�~���^� {U��@�i?���1��e�*8�9tw���� ��d�m�:�u�G�O�.����yM��_�1�Cv�j
�9�m�|��qiІ�t���zc�AKy�1���k~�A�*жc�>��e ��Μꊭf�A��
^���( ���٪�q�\�I|�i�!�*�O}�X��1p0����d���,��E��X�ð�D ��VY2�<�����Y�X�PIAA���@�o9��PH�ҲL���-HA�씧J�8빉�����'��g2��-�p�OX�R�J_֔��m��y�ڧ�	��C��,�iO����hB���&:ǚȗQH|泃�~�}�m�D�9LK����p7V'_N��=�B��׋	�I�7 �	W%س��P(�W��Q�5k�许�<ϒ�I�dbj{?gXͣlh_: �k������%��L��?��\��t&��H���=s�?��0���:N