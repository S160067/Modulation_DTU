��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����0� ����遼�6������"���#�{A���'j�Qj} �}xT	g��F����a��f��洜K%g==�Z���L1������bG����XB�k6T��w+F��3r1#�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv ��i��X��s�-�Q?F�`Y�������� I֏�׋������H[��9����ۍ: ؕ��6ж���Q��" ��y&���Y	6_���.���M�ݟ����k����
۷j	���`a�s�Yot1H���\�뛤tE�v�u�u���ѕ���_ݵo�IF��P�]���=,����1�%��̿����l=���`{逧]�mH��b�����j��Nc$D�xq�Z� �#�S�����Z4�"�o�rF�D�Ɛ:K�I� Q�v ����I���(P�����9��գ����i`�U9@�߳��r\�b0��u&���C�Yd���&P��Af�9�W��6���ak�yr��H��x��	7+ܔ��o�4�
��iT
��*q��-H7��Q�g�ڔ3��o�g��W�$�K�m�� ëG?�
a,/A,�L��=&��h���[�PQ�"��F$�3]���`Z�-�������]G��ibR� ����eU�S��MF����:MiE}4A�' �}�5ΘJ�X�.>L_��v%f��Na����&ӌ'ֆ�u�Z���c���q�0��X���AƵu�}�k�v��6�gIO�~��kZY���2j�n���^�b4�Kݙ�]���f،��D����u�Ű�*<o�3�L
��]��d�NȉK2�F�U �.�ޮ���'�{�#
�1�K�;Ns2����>	��N�&�2�����l~>�� �ـ��~{�����
�~<2��/�+h��X��E������d��G.3�Q5��D!�m� }#�y�fG�g�,���#��]*]q�P�+]��e�Z�De����P�[27j�~�WQs������Pwe	�r��l4��"�RJ�|PL���������
���8�����,�16W�H<d�s�Y�#sF��t#7
gt%R\���.��iX�B��{��	�w�K�v7T�nn����ҭ��MKƿ�/�}���i��'bj �#�{#��'+z}�_⅛p2φ3���fd��A�}�Tkc�64����	u��0��z�6��h;��F;mt8KBq�A?j���2��4�j�w3]����G�֝��f�}3Ї�m��D`���r���k��p_��b@�f��^�h�)-�!�|�^:��yn7)Ɠ���>���ܑ�X��9T<{;&e�|�t��ՑtX!�Xd�f1��i�RK���ɞ��"F��=���V������UI��T��٠76�#��C�����7�3�.�����Q׹���@�>�(Nq��G �\�໎���
P�"WX��3�z���v�zD\f �BjEe�ǘ��cԵ|i܈�X�g���wON�$��;/�9߾�Y��6ݿ�0�����ɵN�x*��w(�ҧ��JO?���(�5�W�����P^ Ȼ��nF"7+�:�s��~T��盀��P�ż�����b�R!��))Y����_Q������e_���S�|M�T�8j ��"ى���Mи�|�[԰x��_�6�1k��MJc�b�_k;��㹍.
9�i�SKX/����s���*'I1�Y�+ح�U��e��ʙ��K<)�d�����F(=�Ѿ�$�)��Δ�2�[�2���<c�8Q1@.Ħ����V4[Z~K�)����ߧ��J���+f,S��y8{%��f����
�����o�z
c2�h",<z*[����Z3"�"3G����uom�s�a#�e=V|(������԰�"p�^���j�Pb
��t#�܌
�t�Mȹ/Uӊ����4���'��jL�UP�q�iߩ�8h �е�5H�1۰y�}�E����r~���Cv�ĮY��z5+&�r��*�*��f���]} C#P-����ob��cժя�b��?��vǹX}G�/J�ﰲ����4y�0���NS'�<;L�~-�B��t�#��f��z�6j�j��J��SVM�g���JmG���-���C�\��.�G;BM5����99��P�l�􂡤�`o��s���atR���Ŧ\Q�k��ó�A��C?1^��� &ӠJ�w�4�1�q����'�Y���}V�5�Rl���މڼ�MBԚ,�u��*�nN��څ/���0��T���}��Ȏ� ��V�6�G���+��m��������o��3׿34VݕB��F��ޥ�Ld3+��o���{-�d�~�O��Q�t���S!?.��#����6Jf��_w�v3w!ɺa����W�N�V��B�TH=��� ��	uN��ÉE���X�=U��hkY��/v��D����5::�WVUt'��b�Jg�c*G]Jn{eݐ�*2�Y�'Y������Ĉ3�m�}J;A�]�I�e���C HBw���aZ�J���|�F��S��1G/���u�5�ƻ$T��Ž�aR*<H��]".���&��m��N�h�:sp�U�B}�PJH������V�*�ȞQ�01e?�7�ȂJ:��t^��s�M�oo��0��qC�%��Ġ��uI�"j ea/�!BZ}�a��.=0? c�����۷�|�o����v�j�N�b&�����T�����;�}X�� �P҆�ΔI�Kǟ�R�$Ƞ���#��\2�{}�=d#�ց�)/YF��G98!h�!V�➷��HkɑsԐ�˜X@N�C�E���'�w��q���rt���w�WO�cp_ T;_-E��nqA��A�k{W�#�s��'	��!�l��rU
����-8{2��P3�ޓ�I�����N9�7�Z��r�Po�}���+�s�3��'��4�]��c]va�)s\8�=��7�RZ=fb`5�6�4U�0vx�-)�+
��������,AASL�u�=�f�w�)�!�5�r<�f��4�Ԯ3��T���Μ��ZYA*�:z)8���2;�0��"�� S�pw���z���lm	W`�����~5(db�1����=��)��B�/���&y|0d��	4�M�h��&�C~�馤�5�lו�����S�T����F����qbl\�[���^��O��Żzduh��)�YUz� ��A.]`��j�*�S[��$Qf�7��>1هA�tt:����\C�>.!�:e��q��W��Fk<��t{��АW]���j�/,q����IZZ���A�nh �����2ҐbhB[Әj���}N<9�N]#���(�QXkk�#m�� �-K���x��ni�$RH��Í,a=��w�ٿ���	����C7��冿4hYH%�C��9���"��D$G��Jd���t>y��x�z��gk,5�I����C��ݚ��?h&eFz�&�~�>l�v�r�(T�#������s&M�2 ����+(���R�d��K���@�73iB㙬]V�rVvd�k��R��Ce]�z�P"��DJ�݉3�i���Jۤ����:���A-�cf�*�j�z����BE�wZP��I��J���k܎!"���ՠ�G%�6.Y�튋2�ushe������|r�������=�8�/5�΂Y�4_ә��T��0ɮ��W�����3��A_��zQ��x�c�ς����e�Î�R�%E����U2����� ��l)׳�8&x����B��`��G��N�Vt�i�;I �����y`���֮����j�}8;��h!A��:�x�}���zi�i*սѿ�zrψ9�.[�M���/�<�43�Z�1(~̦�	��,��~	�}�9��~g`/g���4N+�>��H@p6ܚ�cɈ�)�Y=����Ɇ���+$��0^A����ʬI�F�Β�<�����T�A�4)�-�`U�3��hr>�]-/⽗̄? x�cSE?+q
��]as�����~�]�1��j�)�P�}eخ'�^_��&U�*f��~���!y(��c{���YS�ݺB.�<gP'�N4�KX��n�f8X�@�1��(qc�b��SA~L��R���M�(bh�+d��A���1��E>�#����n/ N��h[���[v���3� z[Iq��1�h�����2����YѾ�{/������h5��5|�K����E[B�K�����Nw�
p�j>�ĳ:g&H{;����g'�v?/��?����E����Qڳ��dѫd���d��~��>�@-��f�D�D��5Y�^�T�_#��~`Z5&`�lO.5�r;jN����)x��F�:4/��"E���-���T���Y��9�����*�&b��晁��$�"���j�G>+nT�{!A�9�,0�WO��0�7��}�M��5��!@�vڰɼ/�����1Iנ�f�ꪻ���,~<��M��D|�6���<mM}j�4";U�[!E�����9a�)���w0���� d٭��2�2i+i�ޙ�N�N���,i���O�a*j1�_j�5�g��3��y��Dl�<n�w	��mPQ���\p7�;���Gs��ݔ�?��y�rO��*�v��~lOz}5�[AwW��]r Y�?��ϣ��iÙ" ���X��ʂ�y�3�YOل���H���������V�A��_-��(��^y�^;~X�Ɛ��7L���<�l�<I<�k{�m��.���kLOx�y�[��$�,"���\�v4|�Ԑ�i(�ݳ����yzA�w�Oi��M�x���Nu��KM!f�U�B��ь��D��s]K�㣂���[�V�T:u=��!	N��EȞ��b�e��eOޯ�C� a��#���cŝ}4Q
J�(/ј�>ϯ}w��w����`�v�����'W+(����!N�{��l�&L87�����Ƿ.��.s�h��������R�6�����}��܅(��X�?��#���,���.�k��k��_�e���a�{��A���͒~�����}���D�p
;�œ�<t����۳oʰ�$*��]�l���߂O2D����Ꭴ�}3�^{#��(�����6&ۄ1�P�%PQ�g*�r�f���o6�c�G�]�p(`]�o$�����;��4!+�o����\��'Ƥ%8HN�\8��r��	Jh��UO��="Ao��p��/]9��X.j��Va�?j�ٿ֑;:1=�,r��9�G�4�X�_г�!��p�hg��~-�1��樌�Y��1>W�,�]i3F�Ԉe�D���F]X�b�2h>��ti��іIbb�_�+L�7���n7�*�k��ʭz��Kf����J�aEW5�K�Mߙ`G���0ܲ�p�=$�Ų��8&����}����9;_���E'�w:֬�Y;���
���uG|���an��J�.�t�5oU�.PX%{X~ql8"�����Y�V�?A@-�h Ώ�@@f��Yt��	k���{��_u��X�n���Z��^�R=S}`7%G��E>#<a���K3R����o	NAPC��?������|R�R'���:'Y���-_�LȸP����u��E�b��i��e���_Ce�z��M]N�I,df���D�W�IP<؀�wZ'�$�a<�r�(!�����jt�,��S�O݋L�_n�3<o���ĳ���a@<t�#)�o&�y�+�T0J��
���Ra|;g�@��ֆ"�EV0z�\�dy�(�����e�S��L�J�4��I�C*p��~Kc���Xj�u�2�K��d"�Kt�&A�Sݤ���/�e�A�\�X{w��bE�l:��r�%L�	x�p��@��6��<�W
J�v�K���XMo�1��M�5a�r�f`zLZ�f;��b��,,DH*=Z��5��>_�W^E�u��ץ��';,��n+c�
�K0MWnni���j��P�5{S\��5�NQ �	���Q�%�n饰N��=����Ñ��M�,�txhb���Oς!�W�f�}���t������Śz�c������n��g�j5?s���nAyUg�W%�|��\�$���F:M��+�߫S����22���=��F�Y�r'��-�M���o9W_>�p�Yu�ُ`�C U��nD���i��#⾹��}�x�����35I�j�y���N7��������^a@
��V��ql�y��xb�`�� �:����|pG���D�n�Ob��e�	!aBl������7�Rm�B��ܯ��IA��&>���hlIR�M�ջ���,'##�<^d
����Ġ����VJK����@�xI6�d��N0�$|��<���N���jC5��������Q)�����<S�z���U\p��Bϳ{Koftx��h�S,H�]X=�icU�2y�e	[/ �-z��J��t�)^Qm�x��ڂ7ûp�����@X58��Ȱ(ڴ����D�	_���ؠ]��ٻފ\���(s�t��_��=�
�p{2���#�Xɢ�3��oO����B-{<���������T����U��U��OFX�����id��>/����l��p[�ZO^;�U!8�h���k����s4�[2i�H�ꬾ�4 N,[��������2_����Ԑ�(���H����ū��1'�JmO���ˉ	�n~T!:5P�!��o��ѩ�9���:��ٻ.LTwP�����٠���_�<�y���/�����+�_��(gR�?�^{�,Q�KSn���C�N���GӞ���(O���=���3��*���Ԝ��B�1�Rz��΂��m:��΃�-��ߤ����x�����5��{�u܀�C�Y}��'}v��qث�M��n�H����97i��v|e�=���,�]�X33���y�rЗk�~z�2r���DP�����(��s<+g�����7e��)���E�⡛������ȠH��\L���y�`�� Q)h�o'�����6TZ�"@�#~�n:�"�q�>���aG��������>B�P�:Ti��� œ�qh�9���G��U)�MA����bΏ���3����Z���_"�}�䰤�ʐR�ｶ�S1(��4�ݟ�9���:(��Y)��|����@	!yG(ts�/�ˎ��垨Nx���u�n�Q�w�]��l�'̫:���q|TR���b-�'E�0:�r�)[؍�e<L�E+� �Dq�S0h~��b��RV��5��z�lXV\ޗT�S	�l�BzD��5�(s����wx�YĹ?��X��4�W%d+o ���e)�����u%u��($�lI ��<����Pou*MGx����/�T�c�s9�AZ{�P!7��aK�Yx�bTy�%uh�o��8�IFN7��+���
Q����eC��S.ܑ9�\�.a����"3H�B��0M�
P�"Rꞑv�ؕ�X��Y19~u0x�c�
$F�f��/`|5�z����.�,b��?���+7hs\ӗ#������Ѓ^-S���c���*���wٙD>^$���i��5���X7�b��b^Gw i	�N�*+]���v�8��kb�������5CA�����TJjh���\�V�Z�0m�Ű
� 1v���N+��<�,D+!�6<Jrߙ'$���Q��@[�H܏'����9�:���1�p���?U��3���ē�_T��R�h�I�io}�
����J5e���0�n����B�����nx�0���!�H���8��^US����&l]9p;E�U�d�>W�#�׬�^�S=M��h %t!O����H*VW� ���(�@����Vɏ�
k�q��Z���h�hs �p{H��)AI��� p+���D�qs���Ȣ>���\r]�lތ�MKB�Q�i����s5���~��ܶ�9�&K(b[��;~%B3��(�ҩ��>�;�%�}���#>s�"�v��;ƻ�P�7�ϘW��6l�+��ךD�.�� �/:�h�=ʘnZ5��8��O�q0�S�VGa7�Eo�A�f'*��7u�b/տ�7�FlY�WeQo�W�����b�bq�J�oe[���§�G 鶒]�C��!,�%I|��JF�G�,��
s�N���8ZB��̎�ĝf�J�'0���68Յg!�L+�+C�
���&�{0Й����Hh��$ٖKC����^�����u^��t���ȡ��;i�3�˄k4je�� ������Ol	���l�q�j�ӛK�#jND�����߿Q�יG�0�JkM;%H�~q�9��P�ۏ�c������}��)}My(E�c���ApO�lh���Aϵ�CD��:i�ۆ]�&@5�˛o�H&��}qf�W�L�	�v���>��ć$��v��w� ^9�;��g�6��?.7�`���P��:����/�!YJm;����~�vk�OGz���	,��.;�i�>���1�-��3�#�v`I&�ɷg����8� ��~>h���t�8��{�P%E�
�p��ᾍ� �Ep�]�=������V�K��\\c�ٜ��-�::�wV%*DD��緵��f0W|(���N�E7[��*�A����y����1����QRVG���-:.�+/�?�o?P��\^�>�dN�C:K��!z� �-��O����S���N��^[��6O�"� ����=���5p�P�^�)9y�qj~�4��rmk��8�RL�Hk A�����F&�014��j+���dj��Q$9�_�e���D�r�y 0�]w��Yi��h̘%,;xg~E�������H䆜�eָ�,��˿�r"���}�]���^���{��!Ǣ�Ud��CQ6p�a/��x`%_�U���L�@�>��Ʃ-H��q��/�@��؎�DŗD	N�Зv�D0D5�8]�[B�b��n�U�4�}��^t�C��t��O�;�]��1sR	t/������hPX�ք�H���x�7��W"�i�F|��U�t�E��l{$βC7�!�H*�琟;���J��G;������\��7ބ���Kal�v��O���lu���nu/t�7bO���#�b��7E����ԇt&�7�����cC=s�B���f�a_0�8OWT�?���\�36������������|���E(P���bv�w���´���fH�\��+l[�`*�3۫JC���W�UaX
���t�^�LU{G c8*�^{(��$_y���fÞ�!�+�a�=��*�]w�*~���5��C��*X'1������*���AB��<ý�#Z	�y���ƌHι�Bn+*q�YM%^�;A��|����+{������L�-E��j
��!ٷEsO�~!��eFo~-	za#�����C�!㕄s4-:�	]o��Q�C�4��2�)�1���s�پ���g:��	��{�B]k���B��K�O�"̇�FC��}��m e�����:��p�u2��F����V��6���+	,����x�9GE�Z�^Ȃ���V�ofC�q�L�Vm�\ݒ�BŪ�|̓�1���)��f�
�*�!w9�n��4.�n���F nGլ�d�k���.(���R'l�ReW�4l�L�Oi4��!�!n��q�&�'��V׮��2����_�T��C�d)�dƲ�
�6%�F��	Eے�X k:�Y��#�-ʬs:w�SF�d�_�С�+�[aR�^�ҥ݆ٓ�r!�I�xS��_>�'$�n	�C뚶ƵT������1�]D�E���o4۞��)��	��$^�;tj��f���R}E��$�,�yI��9w�1B��G��oO��!� w�#�-��h�o�(����M`�����ht��I�V~k?� ��3��@㜡g�eE�`�&P`.�~�?���@cu=�w�K��2UQ�j�/���Ϊ\�kЏ��b���v�*#�[\8_�X�	���Ҽ�'�^�B�R�{)��i��� =��Pݱ��A�;���U��"oA�A��;!�#\B�C&Gg+GڳKu�ОK�	�v a��[@=<M@<�{��U��Fn���➆����n�IZ��)��j� �E���a?i0S;�ν�G̾g˛يܖ>Պ*�����I���-T���wj�ʧW5{t}��`����!�o�&��Po���1�B��m^�J�I��CC�_�5n�]6�5:b�!圖�a��ru��'=���ܦ�c�́��I_(���(�R5c�X#*�Fa�6�:���w'	��%ļ�d��IYg[a\m��:n�15�4��:���-ɛ��\"e�OUo�QV\�:$��*ߡf#¶z��/6}�i�0|(4�d��3��L0���4���He¥�'6Xa����6Oz˵���
{{�Xk�I�i	|�!e�;4OP|��j�����dpy�4�o�L���R��sy�K�����	�{�<���e�Ĥy��p���D�p뜲�5o"�^o�i�d�J��n�`.YU������g���n�Cr�Ғq�x0��Z����1}��˰Y*�n�������8d��QI�eL��8��f �994�5;U���Q�9����f4Tg�'�{�偋R��e�e\�O&"Euv�qSzN�3W^��b��z�ٓ���ٝ�*��5$#M���|�FJ^�����q�J�E����q� ��0��:��q��S����C����us�Hb��@�/2���?��H��_��������hW�8��@�B��Z�4L�c��П�DW
�j�p��J�����+�W 2�����K�f6�����X4&l��\�VyŎ`a�V��r�W�ŁD���z�=�sC+](=gc��Dc�2��:����RH���z�oNx��O�c��7��I@%���*՛��{VEӆ�|�����g{��l���O.H��{`�9B�>��K	�S�_ו�v~*��N��~mSϒ��C}���wV�U��Kї���K.������/x������H�����N%�II��*��<� �"�i�eis��r��Jl`�ْZ����ȿO����B�������xf�=\�ڰ)����vZ䅑�qA^�t�ާ�舔~��^��k�m�hw�M����!��`�- -Z��̍�������S)�k��)ϑ��#mF�GT.�,��e���3~��L��h�P����jӇ�f=?dI��f�Rģ>>�KN\'����1���]�7`����P%�α���E�H�4ⷘ�l������|c�W?�I��^�l
�����f��GF��
V�O�$�V��,��p���y��sG�mU�AP*��cQƚ>�1����~�TJcB��'���n[F��py m�b�[���Jya��}*�@H:h�p��%��2���$ba�6�
�����g@C��t��^h�e��d��� x!��#�S׭������r0�s�+�_(�-k-�X�B~�N�lE�u�n�D3S���`�A+�+bc���X��\�Ap�%�?<'�g��?�v�����Z��⯷�c:/0{=�����U���u��I��ң�{��������ϗ�B<Sb=��"?�=�8��Z�S�b�=t�T�!��2[c:c��pv	)�G͖�.��wy|N�c�/���Z(�nԛxoi�z�2���#|�7���x�*����`�h�S�wg��?+���z�(�h�<�̦Y�� Ф�B�!���t' �Lv�`��\<�})���P�(�n��
^C7��l�T�7���}�0��̮��ʷ��<�ώY�7��O`rM��,�̭�I]��V�DJIΉQ���߾P��9�΂t+ss�I��]-��5���$ou!���DN��}��]�\/i��7�fU��{�<�=�e�q�k��*������z��:uj��N	�,����7�(Js�3aP�<�-V��(�t��zx�*�J#3x��z�z�]���:�����+�����W�{���?@������߭Ӣ}�GP�|ި�V�(���������(��c�4����YI�����7�-�PFw���N24�ϵM`���Ј�Ujx�����o�f0<����4�g�I����W����
4[M�u?�_�l�ʛʵ�G��A�f�Ӈ�w:�Z�Ņ��3pRQ��陨F{�R��{4��~��zl�Ƣ�d��L<wF�&BK��NY_�Cyӡ��o7�`bm�7��3�ȿ*�Wk��7�b��Kg3诒��q"$X+Fb�F3BW���Y)��(8_c�Zh���e���� sĞ�U�(�>g�_-��sW�|UB��{��}��X`k�G�ö	��n�{�'>q?|��\B%i��٤O�D(��ł4U���}��N.���59ʥ��;��Ӊ���BO���U�f�-Ң��������3��Zޖ/�����.o����E�.�)^����I��C�	����6��M��\s|��8Q(����r�',�tS��5�^�����C~k�=�Om��ŝ6�G�xۙ���"�2F�|�=U����:~����3�˸( \^��[Y���G��q��!A��WL��)7���DBs
��K7����Ś�04XA��8�_U�&���T�'�y,�|t����� ��3�MF���r�tQ�8�����|�E�XDٽݓ��䳿!��/��2��i��D �܄�}�<���ܟ��i?��"�M�=���s;B�ؐʦ�8���.��a���i8��%]K�jJN�ݚM��o�d�NL7݊�5u#� ƞ"mnht�{�(�6���KZ�R��э{����շe����VmF���l=\	����~��;#�q�;���f۽ވ����B�ρ^��t��`�vG����^X�.�-�ME	7S�5��6���k�.3��
F��_�wM�8�?�^���8�e����kV�7ʬ��&4��>
��M�x=v�Z��k���+�����������L���	,��fV�،� Ǧyo2��
�T9�},vu:������-��Z���X���2�l�D�"�h(9m+�1E��A��Cs�������{��q7�n�E�@�^Z[l�ԴG���j����! ��9f�6}x�M�u�ʉ�XVO�F [�8��l'b4((��s����;js��w$�9�sy�%�����1AZE�3 & �m�y-��6�"ňEj`���u�:0~+�
���V��g�A�>e��8	ܐ
�e�M��m��n��y"́Q���	�y%d�G0�Ôr���2�dE�ҍ>:���MV|���n��1�g�<�ڐ4�N��Sg���|���N�m�x���/M�`E)���N�QY�r����~A��B���"�݋��J,�C8}ݛb�~ޜ�"�{� Bt�{���c�c�����t�K��$Z�(M���G��i0H�i������Ҙ��_����CU�)�s��Њ.��L�I�az��_�c�����,WJ� �:%(ka��[I�Ml��D��G��ֺ�0+v据��<}���j��<�셑�� �g�&���
l��Z��Z�,^$:��	 ���u�<���y��,���F�e�,�0T'�����R��k��.�y��OZ��pxd����#�����á-�f-�ͨ�)r�RК���E��;(����g��"��bҼ�������Z�3/�f
��h��A���
�:*J�rޝzB������-�h������Ď蟪�8������:*N��J=�S_�����	x�w��êȴ��pkJl柂��9�����@�������=�Gyc� 9�zι���^���1Œ��V�����%���U��V*iD�D�n�9ևjˌI;�EOA�(�����nvZ�*ٮ���u�~<�%>>�Y�!Z;��ۏ�x���vF<ńIP�g0�~���F)�0PG�-�#1�ړ��<��w����&�m�� 1�f0k����,�����/ ����zz3dd'���;d}���0(�Yh���l�<��WI:�k�����ơ�'�<U-�g9�/t�-e�Y��j@U�v�)�xGa�T�C�ύ5���A�ko�S(Ff�O9�\�I��&��,m�ؗiӳ�4�s�L=��k��lZ���&8\F���\�?����,3S,�5�2�h�A �%	��,(��W$(�!�0�x��<]i���K�%N�k�P&��هbK�9���g!�4� x|�@�r�`�u�����e�zX�@����Cc�U�#��*_��!�yŤԡ����A'��TJ����񿍕'�_� x~�kWS.�M�h�8T,q$n~����7h��U�=�%i��y7�]&f +���b r��P��Rdl\_d׺�ڼ��&��'�C��z�@�EX-�Z��3�;�v�c��K�~�_�{�߾��pǒ�Or��͓�	$��nR�k�ۯ�k���.���p��U~F29�3އ~��&[������KA�n�0�ӿ�V�.&�1�b���@z!D��'Uaj�
�~+��|���@f���G�&U�~�J�K�u���l���~k�AD���+�sઠҖo�K痶S�w�.�����>�M[��QC����[�`��P/���;���z��W��֌��J_C�����';�`����4uCٯ�Z���;�6�F��ݔ�csY���U,c��܏U��Z$ϯ�b� @ �DR���(Vc��Ȓ��h�8~�^�Ki:u:�BKɠ��uS���nq�A_��Aݪ�B�p�>�PGo"�o�D�ar#*T��X|��y�q ��W��yd���:�!5:�Uq���7���~�8�<�����a���C{���%fʱ$���_dh+f��"��}�1K��2�$7�pږ�;���A��)8��߷pe�۸E��Lk��?��[�۠�����$���Gh������1�N��4=1��߯cWF�_R��P��[r���{�GL_iq�l����֚[ْ<�WQ���u�I�,���Ij:���
����[b��:�f=Ė�^1My]�'��)A�8m�mL�1��& ���)�jޑ�tE�^�j�gK7�,B�%B:�	}��F`OU���8)%ؿ��f�ŸwKߎS�Q-�B�e��5�ɤM;&�Z4H���mr�U�ߴ����۬Vi�7��o�~"4nb�5�q^�d�/�ap��Z� ߭���M+_�$S�N�
�Ŏ�V��M���ř;%	���tԐQ�К�Lƪ�s�TrO���l�_$��x�/�*X�hS"Qmb1�JZhm���W2��=�0�	�+�R���/�sޒX�q�zh�gg�c�
�	jˏ�GBE��P����O��W�[Ap�ʫM��ђ�^���iM���(9����~���3C�	Q ?#%��qϜ�u�5����b_+��(����]�M��.�b�����s,�%3N�|�^�y���I�-5@�Z-21gZk�/�vFh�#��n�E����}�_S�����Q#Yq��.�����, ���U:�_�ᑛ�n�ݨ=f`�6e�>L��6��&���[*�;�[S���BR��<W�@���c�E<ó������`0w�U�C�C�fXAr3�AR��2+�mT�p��7�1*nk(;e����C{��)U66�}������H�A0;�}���/��O�2��˚�gߴwJ��Ɨs���4{U�V�89���̾��uE]>aH�aqu���l�nQ��}noO�|K�.��Ǘ�q%�	�!��;�5Z.��/��Ҩ�5�Yu����q�(�y>z�_��\P�p���'Pr���������n���X}�*�K�?��L0?�횉������mx���yM抂�wJ~��Db��W����QU�����1r�K��ҕ������4x!U�p$�K_��;`ho�[�s�s'"�D��q�?�<������+�-7`�n��5��g*!����4��?Y�%�-uSX�_��ƪ q���Q�,�Uݧ�\}F66�l��uth�=`��t�W�Cl(��
���B�ذ:&�	r[q�s5�7�`�B�A��+�6f��}Adl09��7?���g�;�8厁���!;5+VS/7�6ۂXJU�抝�_���P����ɩ���� ;�*G��J��&'�q������UO��
t�єZ���Oj���������i{���X��D�v6��, /	��/Q)�������v2���Ir�0sS��O?���F��F��x��v@��J^]�[��6a{J��<���Ǳ`}��*����X-6��"pe��Iu���Nc8l�hy+)=��97�3a!SBa:Co�W�� ���2�$@=�����yAN����*p��� x��':jyd�)^
P?lj����+��KX��@�l�擻5ඹ�Q��0�h-7�%��)v��i��/W5��T���كQ�ҁ��p�?H^�1�se�������~A"f�[0�/������O��.~������F�n�R�@V�5j�4I�P�K=��w�����[%cb���s��m�ZD�ɞ��ë..�(ܔHΓ�W*f�j��ڜ+���4���vfJ�|n�@S���D���G��-Ú{�Ze�������2��H�^�E���W�)��E��;G�P=˫��s�m\7��6J��<#"��eAO����t�;#��{!��X�e褦jƁD��jcD�m4;�-�^c�d�%��ڮ���6�����X�O�na�	1s�M)�q���%�V��x�{k�P>�|��M�cn*{���lit�>�JV�����P�}��T[�@S�&�8LT�f
̋Qn.�Ϧ1ʷ;ϓZe5�s+�M� 4��5�!�.K�~�K4ՙ@�MѢ߻���.s��l��:�fc�+�E,�Q�b�q`��!N��W/�!6ތZa}��^������T��Z�8G��B���B�U����k��ʰ�UW�F��1-"�T�	z�l����.:�<RXmns[t����_��Q��[RU�E���"�3o��$��vpĜ}<�CP-����k(��NH��EQ��d��]�ʊ)�_9�v���Βl��x�؅=m��qB|(Z�"�f���F����Į ��~�8p�]Bh�f}<צ���?һk�]Ck`���&,>���t�zn$�mi���i}⿾�3�c�}C��vz��	��������ާ��Ì�}
��y2��;��촷\�*�6_tI�祜֨��nz��sP9�%"؇;�	$�W�݃W���lC�bY�y���oi��4���AD<��G�� n=@����;S[:�2N������P	D�7s�����SYެ��߽ج%?��`܆�CFR�yÖx�)錼T�2�Ǖ�����ծ)��T����}�:�c��S�/-P̡V�dy�ć?Q^U������ �1�|�dy���RgF�����6őlxO��t&pk��������1U�� *��� �F,KV/1�"�;�Y���à<.��Tm���X����_4�(��a���镮�Ge�`F��d;`?l��E%�����T<��X��S�#��M{���}w��R{8z��̦`t����ొ[y)��.�v��{>������7�`)۫�g��7I�w��#������z���c�k@�P�"����oqZ��[9ܞ�09ct)�>5�~��^��q}��y�;}��fM��,��[LP���1di0;��+ɼV[���Bx����m�F�Y;��!%n�y*'�A@}�+Ei�� ��P)1i�e���|�z%c�3���Jˈ�
�0��Ymw��N�T��S�9[d�%�5�?�a�>�̌z�\�*y=w����QR)}�ZMf�������$���[h�l���n��h�w*f9<G���J>�c�4��1w�������κC��_H��#�jD�iu�+�/ҕ��͊��	�%�G��66��s�4�ָ���A5�d]�ߪ����b�ЍW�x	�W]0�ς�F��e)0��TO��`���[�q������ ����A	T��V��쉐�G�l{���V���T^}'(�
�O��� �0UI������n�(,~5�F2����:�_��	�2�R�y���ü��@�ϭ�UUPj*o���&���|c��354�[����%ez]�{�Y��N�A� 	�Y�B2�¿w��m���}�"��ځ�<�3:x�%/�DZL}
g4�o�����'?,��� �H���>���״���jB��$kڕ�2�)4bo�E��������M7�'pE���\����_D��s��w�����78���S���s������9���C���Sy.^�_C��U"}S�\�5�l!;��DE,�-t��rv�w[iަ�-�:����Z5j%R�k]`4��s\�g8�P�/NĽ�"2�>O���a���ȡ\�_�y7ufr�FvD �{�l��f��CO$x��»�d�1�l|2*�Xd�~�ͫ4 pC�����t�)kԙ_ܝ��j,Y��,_e:�ԩho8�fH�-�C�����k/�����[���W����	�@��~��W��X[���(ha����x{)Y[E�M���!�W ��n-mw��J��Q>𓅱��a��ֳS��1 ;Q�L �(�F��n�A�䋡��կ.f%(�W���U7+GK�b��l���!�蝙�zX�#�~p��s������~��%eK����'0������sƐ4�d��¢VȊ3V��	�ws�`��X�$�܊˱�# [bR�c�J�L��D��^�e���ŧ�F�XA�����8���i'dd���m� HN�GQ�k!�8ਆ�m�n��[d#&�z9�gB]J���D�[���e�I�������=�|G���6�������ڂ^5�5W�4��b'(7N�X���{��>c�0Pm1�������pr<�e^��M:��ٿ�*�c_���U��ͼz�Fm�� p��%��3��HF��ذ��K��` I�	���V�v{:	�ub��u�4��d��$	{a�D)�aL��*�W`�-��d���U��,�3�]�hF�:���<y�y�a�ܾ^�N�Ly'@��i9����6d@��:����.�U�����&/��AN �bx�Ϋ�G(厥�X���K��g; aW��h��}�����ˏ����U;oMt��T�9x���RJ�-is��V�����ٍc�Y�Z�k߷�:�:�*���d���m��{='B��D���i��c����z5�3�$���v�R�Ǌ��������u���S4���^���m�܃����i]���z�i��@mG{1��Z�ĥ[_^j�`Jp�H`J;c<t�Y&��`���+�SB�X��Sx"��Y5@����չdWE�ꦱ9V�|d�10��.e����`6x8�f�dơ�)G�C�m���"ј��Cu��^ݲ� շ���b�}S��_ӫ9dͶ����Vd���9A�Q�U؋�g���ú<�Vo4��Ҝ���H=J��v��O?�QзeP�m�p��i���w��}����'�2k�h��`���>M3'�
���DE����u�S��Zǔ��a!a�$L����M�1�{���ϠN����Ɣ��YT[�&̮�W�4*�6.M?t��)�U�����F���)&8)�� 4�r+�za���v�MV���J���O]����0K��"�w���<2r��y��
H�17Kƭ��E�-�F�7��|�iK�e3�ZړT���f�Z_j4V���C
��#����+����)0C*%$�eK��C[�ֱ����L���[�x��cSL/��D!/YvA�a=>`���7+�J?/�7��;�9�k�/Ⱦ*�!��b��I���-��S#6���.�t�v_������˗_�&&��h0����$n^c�B�hO�	ˠxLX��n�#�{p*���YN��)�2�hu3y����k�/ d���E��.�cJ�'V�ꠒ#&+D�AQ�-;b�ud�3o�-'��O�2׻�\A�'�&G�?�ކX���l�!��o�R�8۹�� �W_)	Sc`Ze�.�����Am�� 	7������I�;�LD)h������h���:f�6��U���J�h�a���r6>WG�2>Si��Ö�g��E��9��T�P��>n�+{C���?�O���l*�W$ُ`0�hhv-�������s1�&��~h����{�[���m����v֜��A�Y��7�о��ʘ��s��!���j�8�T����C��Mo2�p���#b�KȺ<x�-A�:��/x��#�M��|�#ֵ�i.S��)���[X��δ�`�̧��21u��lƌgV�E�S��:�A�pW!po�_��O4a�[������3����s����'�;�\�6���6����@On���ƺ5s� �10X�=DR����w-���hlZ�K�'d����|��Ȓ͹�w�	|Z��x��z�>z�����=}�}��eOQ��1чE�3��E5o����t��xV:�i����3���n���B�����[;6� UBRR�������#�L�^�t�}0�i_�Y�Z�M	��]��!}��*���ؐ�r�C��Q	f�����*��.g�y��y�L>�D��Cӕ��R%��+�5��u��"z���B�,+��J޴C�$�*��o�"%8�Cf4�9�Vz<e��@�'�{p��?���m%KW�@��-�GW�.YK�6�S��/������>��l���
s���ǵ�@�,��F�2����<U�L��^�V�4��L�"��Z1{�pG�.�����Tx�$��L��h�#��|�k[�rkF(���#))h�+�j�q��"�t�[��gQ7Ӫ�W6���ϸ78 i$�����B���r��8���a���hU@L?8
�;�����C#�>�,ʥ�z���wjk#�msDQ A�.L��@�{<="��e������4��x�6��je�l��'�fu��#PH&�@��w��I�w�,J�I�u�KW�q��g��α��ܶ.	�_�zٹȨk9b�?$��G�,#p�m-є��s\.w�H�J�6�]ŝ.unP_QKO*Ef�-%���u(1�R]s�0)Fn�qH��U�\��ab;��8�m�v֎9�1��0�[O�9���z�dY������)T�O��[���p���|r��xѣ��ZnC����xR����m}����lh�L�~Fy��,��3�i �|�n=��4X=�*��P�Eκ�T���B�[�N ;�50<�//��T6)��/�]��8*A������<���0Q�
N��F.D=ꯙ��I)�J
��|�.�0����hmo+�ܟS���l�4�~d�{o�T2:Y��6�^o�`o6�-�Z�βی�̱˺^k�+�k����Q��6B�j����v��=Q�6]����kƲ�p������#��4�<'�%�æ�ǳ�ރ%&% o�����ۏ���4lҨ�Է�RS�Sǋ�a�e�4>E��\8�+�DV�~�b
t=Ae����<���y���IM�k���Xg
��H�YB䇿@�a���;����K�g[�ɹ%�i�A�'����[Xc��0ͯ>Ey4�C���F�g^�v�RLu�ٰ�8���E��;�Y��QSx�x4�ܐ�����c�D'^�����D��U	rJVbjHL�߲��;i�X���K������w�N�ve�F�F�5��7�~�X����"�H`Nxq�su1�|�q:�s�ƽG+w�ODJ�>�#��i.�nXSl��{�O�4���u#Eoz�Ec�	d��
jŘ{���%��$�<bQ�7�5FFp��-s�|υ>xC�G"�$� �: HtEH�("�>U#����!6^tR<��fmL�T]�h*@iЖG�CP�q�[r�ҙ��oC�i����bw@�t��j��d��� /��-�6F;BX��	2;���ց��8��F`���@O
K�|���l��e�q��vf��m@b qK�K�k���h��FT�!1���v�˧��4r�Gj4��
���*��>�pi[���Y�7��/F�Nbj*\�D�MPAav�_ΘK�@��m�2�3��ܻ��WB��h�R�8��O�NK�>���[<5��l� Sq��+�����iP�	
��U��WM�BY̜���z����[�v�<b�AƧ/P�P��v���C��O�9�X5OU�G��[2�ڭ^7��udx����Q0%� oF[r�Vz8�mrX;�� ڠ�D��Ĥ2:1�w��Ů�k��!j�Z���4;<m$����9w�y��a���ҹz ��J�, ����h����W�nY�"�X1�)�����t��./�φ��>�%��1<�γ��d�e�닋����F�ހ�^�%3R&|\.����["���O3M�k��䣈��[���9K�����	4Q{^�v�E+q(�F7R�+5��]a�<�-$�̭