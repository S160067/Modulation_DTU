��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����0� ����遼�6������"���#�{A���'j�Qj} �}xT	g��F����a��f��洜K%g==�Z���L1������bG����XB�k6T��w+F��3r1#�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ�A�O�c9b��2���j�:��HA��?�\/��q�k��#W_�0����J杦�&���£mj��̟鬶�Pf�s5��q�Җh.�k�/��HJGS!]$�y�}�t+��`lJ�g����y;~��ޛl�|TI��_/��U�C��6����ê*�hp\�Q^u�b�B,�{P� G�2�X�J{��鏷�����ݨ���P;c@�3ā��m}r�3X!��;
��L���`�!�ܣ�C�s_��*GǍE��H�y�`
i�o��9f��0�񺔤�͇���M\0/e�z�}�!�Z.�G�$���3K߽9�8#��=FC��>�rf7K�hi%L�'���s��V��5�4Y�=�/�Oȴݱi���}S�� Rd b�'*.8&3veؿ���Ob6
�L��@�{S�,B�U�>kw�/14~KJm�w�.�m-��_�*Ki��yCF�V�C}Ô�	�#2��&�Z	��oV�$��cPq���
����������,��qSq���T�ſJ|����4܇�בP�I��C����L����pe`̓��Q+�~�b��Al�4���n�6���
�b�ZuJ�oX�4i�����sb��gUm�KO�z�-�=4s)���)l0�!�(�������wG��H��v���QX��9�ou䰦k27S��ޟG_�����a�=6�61!Gg�VI)pY|�-��,5�������ºt��Q�h6�D�!v�k\ �4o��/�^�]VU=��V��H�i+��A�vc�@�q�� {d�y5�?�� {uPPR�; ��@E�go��\ 6�~r��%(af$��j�!���>�yT ȝ�h�A�◬�d x�''��8u���Z���IG��� ����������d k��)I�����b����/��0m0�g_9o����Il �X"X��l�D3�KW-荒¥��V$��u���ţ'��(E׹Zh��C�Eī$��
Q@�(D�T]h�8S�$ܕRηj��:��+ᙯa�SP5�,�y;�����I���Xjj����崭i�8ধN�M��s���	A� Yf�L���4k���)�8���6�~p��/.�`���;��_����.y�����"%c�آD	�`�q<A �bL����RK�@�\4�	�:0�xY���^�����Z�l��[��CS/�δ�ߨ@2���
�������y*.���#���U�/'�Y���!���s_Y��$%J?|2�����ް�@@H��0'ZkJNrY3�=�};���z������jH��Ĵ@�|T�ybA�pmb��6ߐ�A���ɅL�ʏ��6�Yt7�,˿XtXTDf�u��q1ɼ��\�g�� f�1��ۍw����U>Pyn���!�b�pe�,ρf���UP��F�俤��-5- V�<��6��3h04�B��<Ei��Ku]S d��+M<,����\�x�`�v�ۏ�8=��x���Ht���2 +W�yG�S�4�͘m���b��H�<a 휮���e���=��S��+լag�sp�D ��T� ��A|Z=�l��|ƺ��*����>��VsεK�����e�� ڰ���{����
QTܖV��;������j�#�5�����*�B(�l"��B q�wL�p�I�y,�hv�_����:o�"L�ˣ����2cT��kgT���4�RD�
���#��+��3�q��v~��B+ӓ��|�=	��>yF+��Ԯ��!���\��'�gE��������jJd�zBq/.�S�f�H${�ԇ�Ǡ���,l���� G���(���O����^�$� 쇎��!�����s�����Lm�\�by��"\@ú���-^�/UR��1O�?����fF�TΑ3�~V�v^��w���#�/ْU�љ���y��6�d��&dw5yVJdps�σ�l[�-b�Ĳ���4F	���^��Yl8�3�6��*���I�1\W��)�@?gaԜ0���K�_UK��M��e����6m��EX�E��c�5�M������Lm^�t�ېJ���ě���RƲ��w�j!c����D��p���A,-6\<��9�2�Ć~�}.�P�$���\��偁s,ˢ2h:H�.2�R{6!>���i��De��h[�9z�J	5��}3�<SG���o�q��zu*��V�k{6�<uٔ{��K4���!��hy�P�8s�TVk�L%��㩪�~D`WL�v}�~o��b��	��������<��	�����z6��78��R ���e�Eݝ�_�󄓇�·�6��Ylw�s��m�u���Gx�)��NmqQ�O�3����U�kv�1_kԥ�_�_x"�Ca����_-&���~�2��_����U��oC�ib�۶����n�"5D���?v�����~&7_',��*G*��p����1;I���H�`�oS���p��H�}�L�b(� +��gpd#o���}��6�����`�EI}wD��6�9]PU���� �%D�0-r`�7j��Z�3'*�{�b�bg��D>�%�85�.�����$�Ι�>M�����@�U��FT�).��ə���k�|�z�Gq����z+$ퟠ��h���d�6I��Q�n��c,�����$ �7?)�r%���C���p��I ��l�7�Wˊ.m�#�؞C�Y{��z9[z���c����y�
A����4�TaW��G��9�0.����鹷�HrE��f?ؘ�r.���b��A�s��W��*G�	��-~������OW�G�d2���h� ��}�mY��u�QsM�@��Ǥ�;GM>�Z�-l���,��U��jE:WNŭ��~V�pG����L�	+�PIPIUCܞҚ������Ĝ��<_��9��U����ҥ����J��di�U��j�࿢��[�+O�Q�X6��9�3����/9�$�� �M�nr�����
���:�e�Ѧї|���Z�����Q����~�4/�=�G��`�
z������MF��1L�d(��e��/rǢA8Ƣ�F���P��R�w�n �vz\B~�N�JC+Lb�b��w�����>FPW���{�y�^	իK������h6�?��	vUW�������G	[�]�վQb&�,��4�W�DU�����G�V]����*f���ї-���[��=13T ��t9PԹ�yH�"�����-��̯��$d2��ƪO}�{2��V@N�=G,�*�N�h�^�%������ȱ��5�Bl��喊!�,;��/��zkg"��%P�؅o����L	'���k�i�'֢��RaX$J_�1N�Id�5jX�z��r5�� �M+� Y��J�ۮ�Os��Fhpj�;K7�\���"��n�xpDry�_}��&��O�kֵoG�g��֔u���`�M��u� �\]{����Y����"6��_�gxt��.���5�Yx~-�;L�1&%
�r���9���ڛcW�^�%�	E�����&gD-B�*��Ͳ>bf�9rӍ!�MO����DҦㄯjT�K� ��목f��%�:� G��@l�<R!�,�T�N�j�8;pλ�~ U�&�0����cQ�ܱ(����ڒ�8�h6��nd�O��hjռ���黫ay���8���)��SA��\�]��6�K}�.�T5���P������䴷Ү�po�@�n �q�n	�w*f���]Xe��]HvK�ֱ�G-�rw8C�s��+��KZ=�ޒ��gTӃLs�����F,sN|/�*��;t�c�D�ݢ G7���Í��sk�h�M4I�8p��r���}��]7�q�)��Zm�޷��I�*p�1J��J�>����[�}x�w���۰�R,fCNdM"�u�@��d0g�iÛ��'�����y	(���c�F�lߺBȝݸ^QS	^# ��\�]�:+���s�ҊUu�Tsđ]�r�}TG�
Q`�fd�LB����]'�����Z�h�ik$� �*��`������Β�{��e>�0����y3e��Z&4��E`��Fyp��On�,Y��e}>jo�C�9���Q�Au�@�f�<�eh[�)���\n�</��J7&Ki���#�]>F�F�:%��?����G'���	1)UF��J���r�Uv;ۑh�LD�S�aD��}A��'�-)�mcyf9��~.�M�v��H���$�\0^|�N;S�==�΁m��c���w��H�X�������($����R�?�jb_�K�n[��[��Z���t(� ��	��������2��5���SLN���6�N���o�=W(B��C�c��ؚ�	@��67̈~���0Zd#�R�F�h���z�Z���aC��ٗ�@�ϳ0���k�%�l`��u�@J=�o��s����j�)x"G8��L�+���Do|�IP$��P�<,絭sE�nj�����"/Ő�O��:���l=��u��9�6��݈�_C��	��dr/��$��h���l1U�3��|b�T�X� �Z�~�I���]q㕤Q��f����E��:�U���X�S%�=�[~�NL_�#geM.T-8im4Z��?/�jJ�#�c<�*���h�d������JJ�/`E	��lr�8���*չ��E���C�����K�e��eRD��G܆���'_�	"����^;��.�a��v%�]��O�^OI�]�^���A����2
fv��\GϜ�%��ta������<IA�|����B2��Ӟ�H���V�g6��1w �-~O��G���e���\���T؝ծ00Ɓ3:Q�������$eS2��:)=��aȳ����H|��X���.����R��h�!_��$<k���P4-f�r-�F;5����4X�u�	}�����6��C;�e��ё�<T��vT���y���B��w�G�Zn�s��3zA�ꂎ �峸؝:�����a�i��ˡ<ݾ+�c�rd������ao�(�?g̝^��O��]����JX^ǕzJO��mƋf|)�(\q��w?�MP�O����i~�~��Ki�)Qs�-DHo�����pV%ܮ���ʚ��K�U�Ew`,t�N�u<m�����<e��~���G�"�����_
��J�����m^(�c�2+N	�r+�~�R��r���1���X{v����� Nb��jc��F���y"W=�ny�`بz�^�?�K93�s��g\��N2����ၞ!AQ3w�z�Gr��݁�����$W�����i�+�d��\���W��h6č�ݮ<�-;���y��VF�VD�t
;F���)�<"vf�Y��˻�����ߧ4a`�].Ԥ-�^�%ϳN?*�	[yH�K��}��4�����\|H9�D@&������K�pl��s/�TγG�O5W���W���Ϲ���d���]V�~��Bm��N���s(f*Ђ"}��wT4��ʁ��l��ŭ�BAnRP��71!��P#����d�IQ��6���
�:)���\�KBYyD\P���!a�ܒ<(�!�l����1Xq�[7��%������W`�t��xG0q�O%�f�lXqq9���`2�>^C�2��{���.�L��:U��r���i�b�G���̞ջ����Ey�"S+u��p�����J�+�%�@$t�"���=�1�O�3{LV|�Ec���!<����,�~_<&/�����a+�{�E�����>v]h������ҭ���Z����a�x���3�w����P��O�M��)6,�6��!�,	~�*#��d�=��+�����䕈&9��d�w�k�(�����}	�o^�O��C��*���ס�G������A��{9�:Dy��F����Y��ݠp3$s��"����]%j�n�k �X�M�;�w�O�z��C���]��r��Җ�J�BlP}�ĦB$8+���AF�$R�c��8u~{W����}��B�HP�-����jA�4E�4�,x_�u�7��zI���*�te3�''|�Zz������L6�eO�̔����Lo�6B�-��
B(�s�y$�|(�;J,;�i�F���/����(֦U�q���*��Tsd����㫋�wDƴ�E@�?�OH�&h��s��Z�ƒ�ɸ������Gs6'H7d�:�'֝'��y�۲�Ý�A$9I��n.�yp)=W����G���k�%�`� �&%ٲ�VȑTFH-?��'\��������ߙ�a�A�u�<�����2a�	
=��Ԧ��r,�^1��r���[_Tƞ׾y-�k0��Vr{�f-݄#@�#��F����Sc�w�7�<zʵ���TR&�[��u!��R�����)�� h���S��ք��1����M���d �&}�b~���,�*��Ȼ�.��Q�񱎜�!�hm��^�w��~����-v8�o"diu�ƃ�;�Ň��A��m�>ZP!x+�;]ty,��m����*�]���uw	��	�TA�'\Э�lQ�����פ���Y�P�+$U=l��,��q�Ŀ����������v�|rlSG���<ꂤ%�����=�Ώ)����AC�����*�肏1�l��/Q ľ6^;�5Y:�����Ī���*��Ԏ)��N<�S�o+�Qt?��gMu�Ho���?spG}q;�ơ_q�"U}'#7vR7��Jq�⶚�o�ʑ�@q*o�p3/����>&�ڏ�R�X�6@�
e������$�?E�����c�árX��OF�%L�{�*y��_��or���z�u�Ҍmh��*����Ֆ��4�}����ю�?3`Ҙ���^�x|)[ں[,�J���&���vE|b%�l�bA��э��'�H�x@I蕞4�#R��G����T��L���q�0�ى�z>�42�&�_~��t�R���![�zr@����S��8��KYb�z���PX��*X�I�Dg'�f��-�@m �_�U���7�c�`�n?
�^�3n��Tad�N�>v�Jc�ޤ���1SOmN`�,oE�p�e^�)����R6���|v���j9]�,Y���x���a�ń�Q�-��[����Qx�����5"�UΜ��1��O��I86��m�?p�@#�U�1g:���6+8+3(B�Y9��[hfhb�Ύ/]ޢppZ���!6&���X��|�߈��s�^b�7�`���2i"8M���H75J�$����+-hsj2���w���cH��������5vj�i��w�˲RUӾ�>����tOĐP��1Wھޞ l�4a]��dWJ/��B)���k�=o�A�u����+s�SL��[ǃ߼y���64#�Fb��i�3D�a�x�sZ�Ҽ�,��|��}��3��,׃K�_c��q��o�"T*9�N#��>o��[���Pֺ�S���|[�6R�]t�KjqT�"$�]S#t񵮮�(��k�ٖ6�g�}q\m�4)}Z4˸����Y���?����}����h��̭j# o�e������t�͢d��I���Qo�Նj����lzplb.������%����B}�����#0��5`��&[\�T;
m�օ�3ҕ Ɉ8V0H׮*���L�0c����sH{�j���Լ��=��.��s���p��o�Lm�?�[�U��=���De�Wp�l��{,C��{uc}��7�?ltr'����f7�<��j1��=��S���Cw0i�2���6�zL�	��
0�N@�2Zl��a�*��K�w[V�X�u�z���YI� &.n�>��ˈ�-�B/�g)��@�o�_K�Z�i��).��5flТ������U��:��."�"�Y)��/Ʉͮ��s���`G��g����-E���m+[�;�P+,
��6� ��0ڽ����t�P7d���D5�&�#'vl�1!2Lm[=��s�+�y����_R���FG� ��߻?V;t@,B9��<�s���rߐc��a�n%�D���u$ق��o�N"-�*�0Z�O�����"a�ѕ�
�=:�����)u�`�'���Ǥ���ɾ���V��zQ=40Z��\�~s����G#F���Rt;rA�Ux��$�yb���Uk��3m�e(���#;�W�G��p���Z{"aMh�O��Md���n��7��ˑ���B4�m��v�Bnz�ߑG�������g-����)7�N�s�FQ����K�1����\�9�e��-��F��,\�3��;c�ܛ�h�J5���f���@��g/�מ=W�p��	B$j��F�:���.Ҧ�3���D#-�I�{O]�9�s��ũ����ac,k��Z�)M��د⠺�r+���~�L�1:Y�U�Ѝ1�^[@t�V���r�հ�K\�Y.>��!�-��à�7zEh����M�/U�*vt5ٙ3�3����v4�W	@�FdP���0�>�`����h�X5�ҳ�!V�N�š������'�$�Uׅ�m�ߩ	��H� �K��@A���N�r=�j��G���G} oM�ޔb"�H�`�] 1u(���`�ɪڎ�g)u�0T ����Q�6�pA�C�n�b�Q�Y��2�������HjD���Ak{�>,����p� ������A�.�Z�m���@?q�;Md���Q��m������̥�;l}�P��Dy@�'V��( $�c���ƻ���^S[�r\�G{��V�y!�~4W
 Q^�pD66_p��\��+��k����|��O|�جJ�ljۘ<� ��b���[�3)A�����u����׹㥫|f¯޷:�r� [���hc&[�[���D�ͩI�w0z�G�?�P��a��d����:T	�u�(a�0A��uذ���fs��}�*}A�6��)�1���t��3jj*Oݳ-�+L�"^c���Uͯ�=P���4Hfɬ$�F���X��L�y��zCL�`'I�Osvſ+���Zh%$XF��f��K�>V��`-A0Y�$~M$+�Q!}��}����G�B.���A&�^<��"m�1	�#��>���<�_`6aUjS��OyTȆ,�-U8����K�cT��8eS`�[֌v�����iW��Xi��I��.Y:C��y���3�������}� ?�T����T�D�9�	)umg��6̡�����N%@��4�9&P�kA=d�a��� �?eMf�`#~�u�[��H��j ˟Q�<m����crH����M�eCz�.W��� �o�`v�'[�K�˺a�UTT�kN+� ��`ʔ�+�����C��p9  e?M{&yu}(��!�l#!0!����:WI��6�����ֽ6sD��\�~�R$Bd�ɰ��p�ۨ�,��μ��ý�!%8���qg�?4�r��E��o��8�DUO�U:�%�F廢�&�Ζr��5�JCFa^ܥ6�'��Y}��7i�O�~'VB�޴!���<�M��s��@)�Ȗ��}�2]��vȒ�"b�?�=F3��/����@\��l�Y*$�	_N�Tե!���@hٍ��F:��՟	��e���׭���Q�ƪ-�]ẇ���%��ĝ�ox���R`�k=�=�j���#/F�t�Y�}���Ü���U��R����R^�RU7������%�ң�I�vS�h�*2���7Xf�i�Q�Ʃ^���`���b�4v
(��(�f�9#�i51��L'�?s�	n8cY�$�XnEp3�Z�J�8]�I�c�<0Q;rPe��ȥ��b�u�P3�}����v}Q�x�)���.��Т im�'�}Q����~-d�fs�m�ÿ�Y���%ĸ���`�WKD��"�.h=�qf�7��킔u�mGDJ�������\�ԝ�u�T�����_���!����T�+&����\_;�U��KSnA8e�q�뷁s�)1�E�~κ�a��?�,?��YvI!nf) ߑ'�����|�49"x��o��i�(9������q�������C6�����?3}�^h$�(���l�y�a$�����
 ���:��UV�r1�Z���|Xi���(��_X��2$00��$L�m.��s7��ⴭ#�H�>��vjj�h�G����.X�׷
�X���_��l�q���;��r����i��?	��յU��il���G�ɒ�<����6����z�]��Phܣ�hʦ*rKK(�r\��>�]l��N�N	����?�w�4�*���I�sK��`� �g�f�e3]Rm7gF���>���f�N/c�����$q�qW���N؂�L@db��h��Ԩ*�=����	*s��ʼ�`�������Ո��|���Q��W_��8�X;��:��j��^kiu*�����Ԣ��Y��@��R��ꏪ�,=B<wZ'?�_M+d�ONNue�M������v�mV�q�y�U�Z��WE8�5�-k�+�[@ϧ���d3���?6�����-Z.J�D�{y&?r�b㴇~d�H U@#㰿��Ĝr��'X��+0g7���g�8�l��q������v�T�d'4G<t/n���`���R5���� ��=ҍ*rТ�]|�kҺ<�Yʔ�`�t$Fk����V�o���f ���&���
(�
�ӉF�~k��Dwl��V�_�ŕ��uŽ����x�Yp�^t>o�%�<P����>.��*�1b��!�2�$f���A.�9�|��N���RIw~}&r�&M�a�q�Y֚�ؾ��Ān�1V���C�M$$�}�t�u�;�^���/��n�Ձ.�Ne2I��Ӂ4�g��������d룚`b|.��'�`$.��d92������tR>��
�}��n5�A3W�ǿ��qrn�4��(������ �C�P�sf~���Ŏq�9�QL%F4���*<B�E8�	���
�{OW�V��G��.��븠P�V._[Ќ����>?�h��:��c챩	������������dZ,�\ςgd߇��٢�F����9K:��3k�dv%�C�$'+�*�kPW$dr���tE&�+I@�ޠ�[��><�