��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����0� ����遼�6������"���#�{A���'j�Qj} �}xT	g��F����a��f��洜K%g==�Z���L1������bG����XB�k6T��w+F��3r1#�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^0�"�|s�@u����[ ����h�A�T(�f<��0���1�fp����י��@����^�j؊P���yf��#���7f5`J��4Iک4M��~ǖ{㰢�p���\�7��P�v}���I8^��c�}YӴ�jg����8�����&`,�N����v^2[7é)Q�N"?��1!�V��[\l����'8�-1��C�5��{聴Zϯ�JjD��B!e��������
���6�eO�꣙m�o���a��D�N9�w�!d@m7�:(t���H�:����'���ȜH�u�/�l����.��m%"� ؚ�L~}k�J�B��h$���_q9���t�;��lm+������P��<�_�?Q�Y�Ws8`��b/�\�s)���oɒ��48�R%��Y�8�g,���1-[i'@�ROD�J����A� �S&�˯){�(QJ�}�x�<�Z:�6���^6�e>N�j�'��~�c�����:�/��"���?D%�qiy:L'֎�#��^_���ͤ�[�ӵ[7v%f,��1���^����q���MՎ�c����x�O�:D���l��u���
9�`�\q5J5p=�B���!��i#�j��
-.��W�ag��0*c��:a{����c��}��yb=�۽'��J3�Z�M��U�[�h	pQ<�� ��dP�<B0jM.Z>}��0�Xx0&����Zt����\�a�b;�Ř-b���J��.M�W`4��R�r��
�y}��F��W�%5s���!�eQ�,���~��v��l5`̾j3q�ˋ��������`������&��_��ӔɣG�E�h�!�P��vC�V,��)�Qx^�0�$�23�3����&��)I��L���=C����d� WZ>.oƩف�0n78����,�	=}� s�r���J�P���j��&^�G��Q�]	s]{���^��ZR NIvq�Í����xe�*��������]٬�T���3^8��_�z��_?Rr�N�lg�kK<�I�/�!1��{	��Q�l4�����ߎ���A��I�УLhG�D0�ҙ��΍,����Q�T��i-�ldC=[��H<=�c�OnOC(���:&|x��i���b�T܆k	z�q����\τ�H�P1�ꔹ��3wF^��
���u��/�l���V����O�XZs���.>���}��&�b3�
O��f[��a[�8����%����Nu�Fn����+Yy%j�j�����lHQ������/�D~�`��"��䔇M��w����d;%"^��F��-��檮y�:�+��xʠ�QU��:a	����"6h�:��hE٥�(�ֱ��W�E��'�V�+^9����#5�0mk*��5-�hS�Y#{��c�l�a	nt(�zq����ޫ��.���n�B��� ���DH�T��$5�J�7�`}|���ִ���F�O4�#�PA�����[��K ��#�ݞ��t/��5}z4��L|�J���J����q��G���̆ZF:��9L Yua�> ��fC����ؤB���,i��*�A�ض��0��q̭8�'3�ٷh����8���s÷=��$%HZI���~[����n���J���
ʯ�Ջ�gcR�푤V�s��d�,�6�)�p3�S� Q�l�U�M�'��*Ƕ>��V$F��u���|r"t��!\��l��z�L� �LA�B���_�a_����E�ڞ�`�V����1��L�Ȭ7��!tD�?�Uӆ�ʞ�Q����?P�%6��_�X�̝?��y����D�Y��.�"5*V"���B��\���F2$
��������	��qZ�ɖ*L�&Ey�hid�+��:jm��K8�੽W���s�v6j]�ÃL&k�:_z�*φD�m[Z={�ރ	�hk�����bFRռ�H!1�b	�o�������!r0w��"jj8�`��͝�I�G�|
��׊e�%�o
�d�ji~�� K

�kT�hP�{A����'E[0�?��Կ-�����>J,1����N��B�j�b!��r������Cɕ/�}�6�F�&�=�v��K=���K��N��3?�ă��
s	�!�����4�g���W�#���D�TR��ݸ�gs�8qg�?�:+�#���~o�N<���|�C�����n�;�ed��=@x�G��� w�kp�G<��VH,�%	t4�Mp�9�
��۔N���A��3�3*�S,�k@h�)��E���J�����t�N�K�rPfaGsίJG�J��8@e�1J�}R��FQ�L��z�V��� �O����;�I�U,��Q�
1�gu�Հɛ7h��Z��%wF:���L̾g��亱�S4����pKx��؈��Q��G6�w@�Ѡ}s\��i���uʝ�����u�l���=�q��*�(�\Q��!6�9����If(�X��!�41�����C��F�� ��e��Ӯ}XͶi�`�?ց���.�Tx���~����<�ĥt�TЭzz_��9R�E���7��� �Z-*l;�����+���/�WP�=����u��?�ðd8?s4���x.%�w�F���D�ia�(� ߷3?D��.,����q~��|cϔ
�pY�Z�[�*�T���bX�8����z��ڴ��wo�q��q}抋"LۜGZ,ZH�Ϧ�B���>J���o1�<���ܕ������3͒�d���3��(��ϻ�$X���:���y���@~���,H{�z1��=����R��F����`�U7��D��oʼf"	g^��lp�`�C jTv�ȿ�$�a=�a_)9ڿ����X������
F"���.� *��H�(K���_qO�ȗ{�PMc��P�Y\��H�"}�+K��E���
���u�B��G��Y�CfV��@�f�K;@�[&���%V�h%��&�����q�mP8�.-�>�~k���Q	
@���?��d:�3��*�7��J&2�x0m�#����u��	Z�����Q��QW�QD��@e%Y�����?ƅCAx�Ա�"�R/}�/!K>bK�{2u�wIjeA�<dC��Y������]O�����^^g���]�;\��Hٯ�JP6;��#k��Y��H�[O&��n:�]��uL��g�`��ΥB��QI!�$"I�kI�8!"��L�#�P'* ���<���c�"��	x�r��4P�+2m'��F6�Q���!>k��=����6�w�_h�� ��H���	-�����p4i���Ӳdy����"슥�D>���v������'��1�j����0����x��b�F�<��-��P��x*�
lu�-l�
��<���JU���]�$݈؝�*�{[�3O]j��_�5K��3;��%H��f�5� ;4�o	TwpF�u=�����Ծ�<'[)ź�"�N�&�[ukFu�� �v���v�
!nu/���/P�*�L��e��'�Q�Ԑ�]��u�Ʈ�0�a�1�3�_*�֥E :4L��q�
JB3
�ܶ�:<�:��7M&�-������ zЎs��E(�K��G�6^�4��ԲY3��*0MZG>�T.4��}����"?����]#��|ae"��5J+���I�6���)��Z�jxP�����L����Q���� 	'w�E��:��-�߅�φ��6��hQ %��l��HzH�\���]�ݱ%����S�F����%D~�Ԋl�k�����\;�H?���YqDJ��B�%��h���ނz���\e"PI�[L�����X���JH�0�<�Z����7��ѻ���ɪ�)ĦG�5[P����_ ���l���y�3�;�3<�2g;OR��$�:��I�&tA�)�I���Su*�`��$�]�;���+OKi�Ih���9iw��KeL=Z�����ιN�d1�W����^�X�+��hB?͉o�����xq��������Y5�p��A�<	�0]ʶz^�@�?������1�ř�>�v����s*�>5�]��J�Ya�p��go��^�L_�X_ �=a�g~���tW������.r&�6!�%^^WM�7����Cc��[�/�g{�%�R��ȹ��N�H{�n����Ǌ@J.sK�s�er�Y�V���6w�H��ó�v�?�	翵4Ŗ	]��|��\�
�W�%��"h��z���m�)N�V���|�NT��B�=S3u�Ԣ�|b��I�`�"�Ķ�8>���e���N�7�zK�J�:\;Y����\LA�:>��(�bx��F��F�����Wf��EXV��=�/F�|-9*!+�S9�큪#ER]q�@_~�JB��,����S�9Lk�f��:�Sm�J��&**(���@��/AfdNt����pc�H�C��6�U̎~�fj-K�5����B�z��˓��WX��b*�0m��Đ,c�tqX/��w�5ڑqB{7�̈ןE�e_d�Z�+�.�^q�A����� �
6eY�l�2
�k�a�PƸG���=WSy�(���j#��|���I�j�[����W�")�m���+�Kuf���{���0�T�rA��c�H��\�c�氭�����jk*�ͦr-�����J?@���G>���0�q"(xl��}�{�oNJ`��,�NR�e¿iu�i�1�(E<yJ@�ɚ�`�\��O#����[�3m���	(z�����H"Pm,�`���eǀW/�uY����G�2�߰9��3E���HW�p��s����.�hhc0"�M��Y�6:����X9�|�ѭZ'\<Ϩjэ�:&|�0����t`L�0	`ek�6e=ѫ{�.B �ڹ/�21/Gv�k$q��r�O����|n�'�{�hO��^6���UHRy^P.Q���VY:��%P������"k`�;a�6L�
9	C�(Y��s_�pb�n���pt�1����$�.3�+<�r.�j��e������[WƐ��  ����z8��W���|P$Vo�,��%��⻺N�K��i�=����f�$F�h6-8�^$����u�5���tY�ߨV ���'lu<�\1W��k	�h&��6��Q9�,�~�Uhvp�=���J3w��0D�nxo,f��Ɍ��)�N�'���ew�R�hAu[p5�"��vw#;B�E�s�7�N>�s�'��=V$�����6��ӧ�L��-X��d�>���a�pдD�f����.\ǃAʰ�'P"&��WM_Q��n�����9砿��z3م$D���������|n�nr��w�(S�D[>����>?J�#ȅ�E��ٿ�"Y�����J?������Ph��^2r��8'&�=T��wyL�(�1b�&]M�O�	.����2&2��O�RZj2���|�|���-ܾ`���Wⷅ	�ft�(�{��`�@�t�5ɑ�㜹[N�Z�� ��r���u�A�}?�7Y�Ca:q��q��HK�۫5�$����|�۸����~pA��(��6����i�G���A��N_QZĵ~�Cϳ�VE׀�1t��b��<�b� 6)0���`��h�o��%f��2~��Ql�_3�<��bO�~x�߿zA�]x�e���G7�����S�3��٨���!�Q��{/.��m��hc��Ai��ˍ�/���8�E_��2��JA����rJ-����OV� ���$z�#��?�yQTU�u�Ǩ�Ѡ0�$tmS�6O�4s�Zκ��Mz*)OGr.�P��R���
^��|��m)l0�80�����@�z"��k�@QD,~6��f�_����ֱ?d�����6Z�$���V����Y�����f��x����`�otm\�ݡ˘������?㞏��;:��uͳ!�����I{z�m��;F�����j5vp3�Mw����gyC��?Tp��䈻�>�$�T�A(�#�1Gώ�'���@����z>:���������������Z}�^%Yaw1*�a!�kEha$���Ѭ��X�`V*99��r߭tR��Nb�P���פ	�
�zHن���=��V<o�Tt�ދ| � ��i^M;vw5Kd(,Pтۚ����KuܢUZn��Q�K{օ���Sŭ���LoSP��g%�E�o���.3��_tjǱ�J��<���Q��+����.�C��� �6�.��-�
L�{�e��:X|�xid����][�RBr���D��W	W��ʸ�_w,q�V���[g�W��Ɲ��KKn޳q58|�q�,i�y����_r�&�Q!_2��Q��
���o�q������}�c��
�[p�����z��H>�l��I�fm	�u�~�RMUMPH}f�����Uԏ�>�_1��V���V�����{�ğ���O��)>*��38��
���0!/kʊ|�~[l��qZ��wzp�5YQƘR�8��ULmh�$�|��� ���n$��_\V��WaN���h��Ig`��V׫�GFN3v�f���PG��^��ȧ�,ڦٙ�������/���X��
�h/��GQ��ֶ*�N���G��d9#� ����N!��Á	��L�~쪳=�\�	�q}���Oj���>�E�`F��ߏ<?%q��@��d.ь�	?�e8}������
)���I����$ZU�V�ڣM=^�����9v���������� Ҥ�L�qğ�ǄʳC�)1Dks�o;a����lr��w@MAήӄ6|�	���B-���8�x)�3�K�NM.�l��&B����Z����J)\&�����9�T��@�Ƿ�w�X��,�$s�ާ]�����p �j�������4�ie�����=��*I��0�yDҢnG�Z������V�mMs�{������(Y��ꝛڶ�&)��8yW�����ҀщG�3�_Z����t���G!�I��y�;K�ieIy��#9�i{��[�j#τ�5�H�-P��Dv��&�*�МjyƏs��7x&�v.-3���u?��D����$���fwcޞ�&?~ �;W����g:��V�����1�7SGs�H���lr� �^h��٦�m�\� �3MC��嫁6ϋG
%g���A�9<�#��|�V�pN�N �*� ��ab�'�5����&��m�n�\G��G+�o�Z?�u^�WK��%/�֙�涟Eu�t$��ߛ�B��"yKT�HT����54�|��(�{���Z��W�#͈��>�sZ����I�}x��J��|��E�m_Ӡ��gD�bU��DV9����Hk����y'��>����\Xn��TQ���)]�Pp]��W�jM悠��Rߪ?�eEr����P��N�?1Du��xr(��=DlZ���Gʃ�fA4��eI�H@>(>�I��_���9Q��P�;{j�ɠ6U�(��Xo\��I�ba�[�0���x��~D:����|����#͘��~W���3�ĸBѕ����A�&C���^oG.�z/:�y��T2fp�:��c6]��ؔ�
�b�l�@��i�g��WW5����(N�قF�	Nn��4�4�6�k�D7;ף��*��n�Ƥ��I���l�8�8�b,S&VK�d��܈pu���:���9�»��� 	�
�k��y��)�a��+7Z�Va��L���2�y�,ſ��B�=c����!@@L*�Rƪ:�:v���ǖ�.�M���DJ>=����@�S2��^���u5��蔲G����f(R�D�s��f/��C�gYț���R[0Ggh:�^�1�����\Q��e��X��Ā�B(�@��e������j"!�<�g$[]#��5������L��lby3-���%}�� ���D��QB_�r���_�z+����Hx����]S�=uyx_B��%c^�L�JF�@깜��(Q�����{���a����j1�����-��b���w���h !���i��%�;��	;�(��pհ���p%3ޜA�C��ztU���s���T!@)�S������ໍ]+�m�����`�qyc�� �V0&!��F�3�j.jznR*V�t�QGe+�7?!f{�u�Ӵ�ՠ��pgjD�ʝ�u>��lB�pL�.������(.gk�g׵1��]kص�]ǔ��$���'Px���B�}a5\�r
P�(xX��p�~i�����,��+9�a�G!��U���ݷ˗�楠����B;�E(�Ĕa�"�����	�o�9g$��S�k%.��E���2>����+���mzz 41�z,��;pct�v�%�N9~�կdcH1 ���y�ȌT�s�"�YmO�L��v��67TR��N��k�*���A��N�hS,��yWz����p~����b��^�آ[�t(٦�k����×��j��án�)�����]����!�Ku��z%ݨ �Y�l@9����@�2Й���qM�:n�-��MM ����0i�(���l-Ь����2NQ�y�����RB|1����l� ֫1L���qp�5J$��(�4V�15����ꢄ�R�����r��S���9�q'w���1pBE�C!+{a�3���������+A�P�C�O����Eͦ�q��y����A�U���+�9O$���p���|�hNq��K��ָ����T��E�]�m��ȶ�l,!-Თ%t׍����QN6�gm����n_},3t�"ٱ�p1D���"K��FВ���e�q�'��ҡ!8�;����{JU[�]�Qr.��x�STKu-�\�3֢'�V����܉�;�*�����@36y�霨vf�x�h�i]શ�[�Y�{o-m�>��|�D�
�5P_}ZgL�(Y ��j$��� ��\�՘4C�+����k�6�.L>��ު<�����:�������+�VH���w��E�� �˃��V.T��%�K]b��O<����o{j�СK ����ۍ���_	�I�S��ꦆ��K�kt9ɷ����޳��Jò��kWy��b�\�&��5p��y]H_$���s��D�2�����"I�!����r.y�Ɛ�.MaO���a��2���u��n�-�&1x�t�Ĺ�^�	�a�� ��g��t0E.&�ðB/��E!�9j�%?���Ex}Ub��Ɖ;P�;Dw����:;F�4��p�T�OaM�g��C©���W��,,&���܇#L[1���v,s�W�a�����6hk�[�w�{%�������JV;����i�8��o$�a��2]��;��qh�I��"�9�´��QA�V,bR��O�f��B�i�A����
6^P���Y^���ȳ}��oGe�x�A+>��0MZ�DsD2~�,F�u�3�ݯ<uD�9��)ԅ������-�k�7��*���!F��e�!0[*����΃70�X��9a�Ҽ���O`�>}�B��ݓ���0v)��i	�qq�c1�C�^�e�j�-*ߐ��IQ+Ms�5�S�W�;����4����~���TO  <�i���%�5+��>䧤/��;�� �qI�Yix=q\��!�	���כD	w�x5A��&���Q(�άi1\<iis���p�H�ThJ��M�O�g���&�гΜ�� 󧩺�@�LӠ%�/]w���?�4�1�����u�Q�la��1���l��i�79��}��rg�̀ƌ�(��G�4�(&��W�L0{Da��x����� �Dv���T#�n�-�3�!+�c�=D�+�A�/�J� g����v�mKW�8՟$��f�Hv`���#C.<-�>��p�- #�p�u�}�|��b��S��6��`o�+��,�#N������\��n�Yd&7J;��Xh"2H�%UcU�w�.O^wm�:$�����b:D��<�f��wSy5���[��8���t���Wo��p�j%�:��)��T'���|RGO�q'�NQw�WLG;��������FI d!����_}<)���%�K��0�tkW���ǿ8c~��V��{�@@�z�f�,@��A�Ԝk٦�Y��9|3a����&���7e�!�-éY��Wf;ɍ��:Ι%3o�Xs+uE��e�Z3����Gt��3`�
~��==>G��G��K\��J�d1�霵����|O6`���z�Yv��:Z���䛢8���|���rז���\���bo�'��10��	gЊp�7&IГ0\\�8�#�+��)�|t���n������\lF��z+ڛ�N5���W�m7-$a�����ά�)ǥP[>�&'Uv�a��IQ�3�\����M��ͨ���Z&�D�L�����GaK��kWFĹ~jSvJ��[��5p�QXmh\u��	�]
���l�Hwk�n13��}�n�%s|��]P�Jx�����ԂYJL{z���׏$5���`�Sm��yyo����M��`��}�[��C*���E����Aq/̠ƙ��	�ڛ�I�P�[���r����p���:����+p��G��Ĝ�HD��@ x��B�N�^2%��=��Xd���O�S�ӌ����N�N�jף�,tsꈀq7Yog���k�_�y/+u���"�-�g��0�r)aGp��%�E��?I��;J&��?�gw:w�=��T1w��E��]3��>��JWi��z�Q^�K?���M{ �I�a/�m�9�Co[i��ܶ*ź(�'�Y�%B�C�X97�E��dR9b�#>9DJ������s�0�*2�vR��xzs��|���P�e�M��` K����DN$����n� ��q���;	��C��3l��d��qx�����8̣.�?�����f�#�
O�IP��75/G �*x����UK�+�op.�sC!�\�����:��A��v��Y,��Ɇ��"Q6����b 1�I�{
@���E3
�Au��kl�$���DXޝd�GHQ�<}GaM��<N��ͅ�!gZ��O�C�,����<�M�X�++x��d�'�z��t�ĨM"L�pLξ7�?�n$Y/&�ӯ��.���[��q<�җ��jH8\vhV�}M�e�_E�b��RF�j��a�$F��J.�co̊˄)�G�ҩ���n��X|��;��S�|�wϥ�)�ݓK�� ��\�� 3Kk������{w�"����Zz�� Q�YQ?�(z3�M��־u��(ҥ�HxJ��/vʅ�H������U>�n�G�6�3G��.��=��぀�mr¥��:`����=��e�:���M�_<�KL��|�F�i�!�����R�:���2�t���3�ƚ��SԖ��0��P���@ǦB>m����Y�����jk������apw�����+9�uw�v-^��!��dI�m(	���Y[�X8�䙺�,]�r����7K�.�d���K�u���w/����著j�Ď^��+�3®9ʉ�ԥ��v��_l(�o�����Ve�����\�OZL<P����ٟwB�	��ǭt<�W�Wy��(ĥ5Y��u �$�ҟjB�����ۉ@�����xb ���։��g��~at,
���Wy"s��U�lz����ﰉ�ِ�
�!�j����M�)x�����w^�e�S3$V�eM��� ���i-�x�Jh��U���eW�R�Ua�΅�2RAyx'�7q�m1�V�
f@y�� �1Δ��ū�	���ߟ-V��2:e���2����OO?ƨw���漸IEG�!�֧�u��j�.�!�N�E��@�4������p/m��ڛ"H�ݸ�P1I5K짟K������_���S���Z���%�8@���X���!����v���zj��<Te�t3 �BY���v�D�(���p9?�52݊��Z"�f9�k*a��M�]^Q��Tr���Fn�d�+��é-�Ң	���ׇ�c��I�bC@��bt�P�ބŷ�mʣ�Vպ�j��.s�L��2���:������i��	�Ӣڜ�Ձ�z�U8lPr��0:�u�H	!��?�;�
�����IPdw�,3�jtsU�t�85NL豬ߚ�4oL����,Q��"�Ē���q����^-��z�^���4?�;D���I��A���75����s���8䒢�9�i��\�0������+����L�S���Ir~g�S��l�Pd�M�1�x�͸��!����>���'O< �����鮷�G���Eq�y%��$>zY����|c
Fz��<>�;��b��v:��ؘ��j7��6�p�����R�4`}؊O����T�W4[�j�IC'�b#������4�O�?�u��|'�S���!mf���]�Am���<2�͍�Ѵ�]4'�d��{	(�$��{����M�+Iq�xmN�[�Fa;B�6���1��eڤ��i�<FoQpa�>ẞTz�Ѹ,q����=��P#�aEL��������4��t�*�]��Y��j�''ɳ��!�	���s�@���Z����u�@9ԱN�6�k���7U��7LkF;|�?�)Q��)�-�a	�*P���^ةY���>�p� �V,��L��;e�7��͑�\���&���k�⦱O��HS�}vG�pjKv����ht[�q/���,E^������r�	�;�)m�Xl[�؉��;j�h�����ݐ�ZW�'p�ȟ_{��3MS�����0D#��zH	��V��ZI�
)Ȁ�K�����&`���?]���S�ƙ�u���MY	�;�%Gn��4�Q�:��Ǜ���? �W�*�R�<�5��38``L�ϑr1*HS�*g�=5��gU�Q�v����b�r��LKn�Bn�D�w�k�"�v>�&s�1<�h(	=4�*_��Lh<���I�J8�t9�,Kk���2ߘ7��h���ï>��`hw� ƞ]�(�M6���n�N%<�>R�cqT�5	�㣻��E��r����L9�7�&�q�?A��Zt!BL�����s��y�/LBn��b�3o�2��򄚰y�
�2�Ю3���.��W� ��<����&l ����4[��p�E��YX�)�9~C4��P3*Y�/9�m�,��	'����Y��B��nc&oѱ���2��G�v���2�u�Kl"� �9-���,�V��誙lj��^�����ё���^5��7*���̤Q�~E�N�v��w�#ܔgAT@��Mi�	u�N�Ĺ������nO�=g�}������~C��Ң��`��-?`��o��F-����e˃�" �<]?�NذrA�hСΛ��)])b�b����ɺk�7�1T"s/jA�Ȉ�M������(遷��D��Z;�@�[~��G �����0��Ґ�ޑG�az;� �x)u	+i8�=�a�M�Y�!m-~}�6���%�!�MD}((~8��fQ�'��>NnޯYm���(�Ԭ5���m|:L	��)�ߜ�E�(2!2���g�b�@͊R�ߦDe3{���z���7����7R�����P������j%�&���aJ��%/���8��9��a/�+�Ўm��K)?��[kj\"ݕ��'��©�	�w����5`����%T����k�Ʀ�,tF`��䡃>��>��M$�mE���M�l�h�{9T�(CwJ�z	wL� 0	)��Vݯ�x�/*ϒ5��ڠz<�*L�%��~��fQ��!���ēTm/Љ�9��F�}6��zr �'!���J�n$�RH�,��6$eK���6D���KP��l^J� ����Li��&q7����\�Z�43���C�,��ܮ��$�^Q==���ݼƬ�C2�����RΌ����r���j��w"��@U�5���m�&�B�u�0*8�S>	����%��7Â�����%�)����4��dJ{���HǾ3_���bJW~'�h�+7$�`-i�c5-�]�4�]	�E�3�4�D�(��E�Q\da��9��L-#5��Ʀ�x�T{v�uZ��X�B��NO�Y�#�z3���c�v��=��t>���iP�ᶑ�� �J� ��"�@�H?_	�]r~���/�#��\FѬ��0�w,� du �u<�dbo[[���C����=dd@�g���f�J8J�Gϴ��{K	��<�1V��!�S����x��}���ҏ#eVU��A2I�����(����-|�.B|<ǀm��wp?��G����w���8	E#lh����)}SX
�,A�@�a�5�>����{���ku�5���΂�C��ܝJxt�(|��c��|O[�i�/���B|&��<��%,�u��rm'Nb��i�!�����������=X�"�֘�z�!1�����[Jg�v8K�H�e+�,B�3����Y[�2�&e�����2`�z��S���L����S�%�ǥ~��NC�mE��_���R��-
ɨJ�xg�"l�dԚ��y��p�&�?�>��E���cg�� ��<'��$��ջ��e�^D&�yE�%�~���n
��/sыT�m���0L/�r˲=�mgx6��#�Y�l�$���F����`ԽQw�	�H׏5i����B��������h��?X�	����l�����R�y�N1�l���A����uxNq�/�No�@U�>2rŒ�*�8I[���[�U��;c[�5��2@�S���xw	c�4��O��I2�8�(2����J�ed��7��ʸ^,�B/��k�9��x��n3�_�Ը�!�
�O��+����$�'2Ҫ��UK�ӝ��t�EX��k
O �˺ȵ��Uo�'YV]�>�Z��	�kI'�*�~�99B�]穃ؿM���g|b��ZWG�v��"MxsPA��84�PZ��T`��~n��=�5n�����b	QS��*VWKv>�E7 ���Oi=�o2����"�xK�a�/S�a�a��j3�h��dn�u@�	ц1jƲ{5q�Fjd�w�	�����*L;Ώ��Xŝ�Qq|um������(՛`��Q��T �ߦ�B��7_KH�y���}��X�0P�\̓�G2g1]-�;�b�e�W��I�&/�W#�T6��v��k1�'�aH���V�[�fH`�bmA�QI�Ȏ��y6t��e���mQ�Hο�FFT��w�9���Q�t�c�?��P�OcC�&��A�~�I��R5s���������&���Թ
f���8�:�0U����/$!����>mt�ՌC�>&���m«�tQ�<=����mɡA�������^�� (�7T%�g
��Qben�U���?�^?�*�惿�X��YN�Ҧ��J]H\��>�,@�U�	��	�^��`�o�r:�ߵ���	Mu��$J����V���Yl���I���<����"�kGw��hS���%��W\�B_���{����!K)�357��x�ф��h���I���tW$���h��vʝf �?{<��?v6<�u$ �GL����\�M�8�ܗ�Dg��������Y#�&As�f�ST}=/��5��6-f�k��c�,.�=��Y�;�e��ɯ�0�����Ƴc@E���M�v4����E�\���p��'�ck|�*���W���ã��S���v�ӷf ������f��`>@�i�A=U�!H!�f��"xk���?0
I�1����������w�W�m����������Yի��2�C��é�8ڢ��p���i�$�9|�P���5�>t�	���D��F����'o����-\BIX�mx��3TiU2��N�k�Q���Rz�}~q�+.׾�rQ��K������Ϡ*�i�[A-�y����tIV*�2��ę�?�N�����ĕ��J�������.��:`�y�\�(��o�Q�'����d�G]�ѧ�E��Dr��@[�ܝG����v"urC(�]WF�kP �R4��e�{�0��[������=҈��˾�r���`/l6�z�O�j[Mխ���C�ۗ�y=��n���H��I�����_M3S#ͼ7��@�B�m�|3T�퐶ۜc��Hf&p�Au-q}��*t�x��cŏn�Lmh�20.���-I{�31�mN) 0T��]'�j9ύF�l�oM;ȷ�0�L��Ա����u<��͑��W>Vݦ�}�?�h�&�sNN�3���>��Y.�>WsO��+	P��Y��B�l`F\�Ej��e0i���
)�%�vڿӸ:q�8[aj����[v�c00���h$�h�plTv�f�t�u��&yq�vb0d�D��Ȱox�	R�h���(Q���v_>wfI�'2 �U�,	)��1�WHq���;�/��-��	�������@�	qxO�۴�P1�Ged��v�8��f�!��8�1Q����|Х�X�{������d ��u��"�H[v�7��.�>��Ѩ:�1d'+O;H��K�iXt�뤞�L�i.�H>�\oJ��*��A¿T��%Я�}>��3��l���]o�[tO{�cY8A'�Z�ѕ���h���~F8�t��?�e�Жy$�u�H�& }������c#w�`{���fE�V�!�J�I���%�1i�G!8�G��#�]�dx�r�y}�dt�$� �0X��
ܢc�T�bJ�E�Ė�5��"���"�'E��nw%������[����h�~�p����ጎ|W<�'AY�8V��x��(�T	K���������8Bd����j��=�	/�N�r�׻`հ\?���*	&�DԠ��e�57�Y���O�?���r�H4����ܰ�#��kQ��彦����!��c$: �Tՠ���vӌ�z�D��9���jER���(���SL�u����/��m�`eT2O�N����VGS ���}y�)�&�-�&?kC�^�+���O�+�.�05��dj��M�$��@�K����*��kb6ߌnQ���!�۶n�e>�,]o�W��qM�DG�
yKh���x�����rH�j�%J-E%�6�X��� |�̪A�z�s�8~Z������VlGy�=�7S�$�X6(f�'j=�� ��~�8(7O�5LD ]�Uu�t�F�L> �q�q�ٲ�U�+G�؅:�X�%�T�˸�[a���T\:���9����N�=�V��J�8u��S�	ݘsD�fj��XO�h�Ƚ�za�lNH��F�3\/��U\��2��M؅��3co8��*�yҎ}3�
���9��̭13]߄���M?٤~�Ga�%ͻ�����l��9�8g�W�Y����3������Lz�%d�x�B��p+=7��RlKK i�9���Ѝ�"A��Z��^W�y|��4[���z@	!5���2�J�l�g��dD|B\��g�c�'�C��N��|��]O�&j��Q_�i~t�k�,*����L$���΍����}O w��h����(ez'u��_�3��3`"v㴺�<V_g�F[VQx���մ�Ⱖ�3�TX{��ZG��,\2ƿ��5h�q	ro_h �KJӹJ�(�C��@{�X�_U��1�{�d�R|��T�`r%����s���9�>j�r:�?��w0�)��ϭ��r���)��-�����;Ҧ.����GY w_�AN�H��CdX�c{��I!��i��!,�g˷��K��\F�=2򀝏y+�F~ɥ�N"�<�#��+VǄreAХ4w�]��ܚH1Y�E���P�uy��=1����Č*�y��yR�IpS:?&Gv���PF��3����!}��p���h�SI���s���z�^��V|=R�X����pdQm�-����s@{��h�� �y�b�8�Q�����.���%�D���ڳ�e'���'|���G�źX�|��q¤�!*L�0����:����\����'sD%��4ݗ��|���F�=|��8伧����R�W\�8��G�H��7�{��?L�U[�Z�y}|q�31W��R��fR�\�~��v��|�G1�b�>�k���Ou?��/4}Rwܾ{����!;�p����",<K����iz�0��w�����Bxo��r������B�o) ɭ1���5�Y����2*��J��;�3>-��3Wn&gRً$�T3�b΁��@7Z 8����*�D_.G⍶p��4���Р؞�����;��K���n��a\�.����8~����R?Y�~�ݹh+����Np���)���������jYN����sj-�X���Rd�W�Yk�Na���m�Y�9�ᯪ�/��r�'�kB{��8Łr@*�d"�T���Um�ҙ��{�5��F�xWV	ݐ��Y�r��I���L`�v��2a�<?T�0�e-�CQ���k�Q�y�Sq��~.=�`�_#�^��
�'`\�&�����y��y�v◱�T5X���$C��D��Iߴ[ٜp���%�IdJfjD�{�x�>$��d.0��2��1{�0
�^ap��}zJ%�j��=�h�LK���2:�퉰e;_=�*��9�4����`�59@j�e��K��E�3�Q��v��Ƨs�g���ڠY��ca�ݹ�:�6�Ce��]�s� ����2�h�v��������Ӷ���F0l�eȦ,_�'-Ы�ҧ">|��0���`)gj��EV���y׸{�x_V�5�T���VKA�=1M�sEɸv{y֑>H��C�y�w�J��C]�ȴ�g3{�<$	;m��g� P���P���L���^-g��ЀkJ�P���P���M"�ж��h�$r�$�"�4�'bZ��+Ѫ�>��H�S�1�(�>P�9����kw3�{��|��Qϙ�ۅ�Zݲ�J��c)^,����e�^��F�p���K�Y�]�r$uwn�x�Z���4�#�kR���O!�U( �^����!
2�l��ˁ��I��!�$�C�ę�`����O�l�`LX��J�xs�46fT���%6�諧�K���e�3ĿQ�2�Z4��3�l���+��5"фG1+gc&��|�ٸO4&������B��g���擽�����v�3!��Em������S��.@��U	G{��%_$Ⱥ��xOI��u_�Ge|����Ԉw�㒂I;������TN1J���� �)�pmR��]�=���������>{*���솕I���=�y9=Rm!�SL�3���x��o@VR�1A�s�>xe���%1��_T�� �`�ڎF���Y���u��Qΰ��	��5��*j���<��)
"Mm)5����ٝˍ4���dW�W����ic�b3���r�6�D%�K��`ctB�Z_=L20z��k������շ�1��@��H욉;/$�3,*��O�=^T���ܫ���0�N"���fBΰ$�`u�]\�UbM�v�`�J8}�>��,$�	(���֮&�0?߯���"U8(�bt�Ɲ�N�᭬���P��|���@�p�6gֻ�Nn;a��-�����'J$^�6���Y�2��R�߆G��3f���S���O|D��Y����r�Q'EZOaC�nx��=�|�3�=}�=���#h��Or��*������WRi�D�x�l�cB}Y$�~l��/���� )*�ث�fYa~�.tˆ�/�T����U) ��9��:�U�ң
����F��eC���R�2Ӎ?l�����;���柧��0ks̊��ɤD��9��?��F�
p�'N�,�����ʚ�ބ5�刑`��V~�+#����$b��@~=0{��{W����㳛����S��l7J��y�x�;�����`4=��8@��2�;!�Cb3������t�Q�*��8����v�Œ���m&��4r"Qn�|�[�e��-Y�h��wqE�U�o�86w�ˢ7�b��Y��OZ�O�h���lU�B��JĢa��A�bz_������ $���YW�+�MO��)ǁJvz�b��<l'c��X�"h��v�ł����N�xc�S��n�oy��u���@���O�H�E�����=w��]�l���'�W�,huE�����/�R���S��K��;���ޛ95�����TG�xdM��ǜ����9�CH���3