��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����0� ����遼�6������"���#�{A���'j�Qj} �}xT	g��F����a��f��洜K%g==�Z���L1������bG����XB�k6T��w+F��3r1#�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�A���0>�kz��/ �_M��<-�[a�%�����'(�S��jS_�,��8��T�.B߫C|��N�(ݝ_l0fS!��mYԥQ��DF�S;���h/��9mϓo��ޗ��0���v���(����"�6�6��Z���/�^g�)��<���(�Bk�M9EV#����f��
P6�f�W����t�VF�Idh��,��X9�Rx����������S�.Y#t����WztK�L^�a��S�/[�y������#ғ.���4��'B����Vv��u�$]qti�ԗ4�:�dy�!�&�`�"$pC�V�R��/��j��ч��=5T=�̭r��;���I�vJ2�XaF�-� D��#8�����
)�P�|?���b�+��G/I'�@@���ɮ7�	�O
������nݤ�S5��/�k) ��}�N9��DI_X�N�dՋ���>_]��(6ػB.m���vIz��ͺ*\8v�h�5˾���&��o�a��#��Qm��m[�:��>=�\����Mt���0�9~0����{����� :m�?4!�",�RgmP�9��?9=Ӽ��Tt
��&�RBRq�Gf�@KM��k�Y��4�&M�MO8�H���.qwO�����{7��#��v2���yŦ�k�S��q���x�]�A!���Ձ��ʭ�$�y��eW��f��r�i��zVC���ѝjCxY�V��.�ͩ/�Q���3Y�?`P��|Z�6J��CK�fj�N-ju�=,*���WjN���<6��l��H"��~&Щ_��N�ņ���F��.�H&���>�f�VF��r����m3��c�'�'�9���ϡ�������q��ü�h�B$�+���\1��Ct'���ٿsϤ��#�i�%B#��o�Lrp�����F��:ǖ��s�N*���=<˭���b����ߗ�e�X6<14�t�4��v:m�j )1gH�:g�
'��qʹI�iVӠ@l�m����\��<���;�J�!#ҧ�.-�e��L�Sڏ����_�}�>��:��j���ۛ^��NU�C�b9wzm�|KtGu� L�a}m���Q�ߘ#$�3����ز�Rz��6j%F5�}�V���裕fcShl�c�ի*P��.�c�I��U�Z��%�2����3�tJr����ڛ���zh��ڛ?Yz��TV��d8��� ��K4�"H!���:�O5���"p�������{�8��k�������864��܁�筑��Tpdv� � ���5"v��Q*w\WM��K�$c��%���-���V��ͨi�!�f�o���w����$|�ٰ�a���mb�¥h��^k_U*�C����:-Rl�����=I������I��S���<ꕎ��R	 ����."X�^'ܽ�牕?��u���.�"�T����4 
W��=.�J³���b�8��,��R���Rzw����[ ����ܬ�0����C®eu��C��@��V5^���D�Ӭ�������{>�?�q�/����A8ns���L�ؘ�nSN��Já��a��
�}%%��-^b%�^�/�-���z�ֿ|E��B��w�0���ާ���j�a��h�h=� �Cds����9ב"F�FcW!~��A�nl�����q^7pBB�8ne�/�w�D�t����f>�)n�3�W��#p��-*��[t8{`݂3�]xqJ��"�h���I��l��tYd��RR�@0{�q�o�%��[�l���O%�"�u���_FH[�P޸���I�2ù��V�@�ȣ<�K��OUpE�É���X�G��{*7�J���T��fz$r���<q���X��'����r��{��z����7KB:�� �Ov�so�RE���"*˵]:�A��ɻ������m#s�E�iXQ�ٻp'40�ڦ��Mh/����@ã��[��Q��kz���\��ZR)���xg�%�v�W�ϣ���fxO�KZ<��+�De3c�:'��{u}���H[1��}��/�Ez�)�zW���n�p��0�fe��q-�3@r8EZ It�9+���Qz&��ɮ2��e����d,��$�Enx}�ipDZ���;D��e�;+uJ�D�����(B�����<�a_L�p�N��y.�T64�47|��0��:*�D�1�_.�)�ǎ7!l�F[�| ]��=�i���G�������omU�,�_v�d���9��x���0%R�[\u�sq�a���|��R������Y�6�I\���P��۶(;Þ�ogҞ3���=K��7������.�Fu��f&]M=;�YK�e� m�E5ۡ�H�X\�PQ�7c�3@�;��v���Z)~*z�ʄ�H��4>%o.��8��:!Ͽ���j�}�������ʣLK�_C"��W��~�`"J�ʥ�h������u+J��J�qb�U��p�r}�&-�EJ(j�x������')���%�hY�9°�O�z��E��:z�����V���y��x�����$6���� :��\5,����UO��}�wh�+[����nJ�9$�YT�W,�wl&H:�q���'O3wwϨ��OdAmN2�[���,��P5�gu�χ�F�����S1ֱݬD�_�=D_��*��s�������\'-#Yf�ZL��	��|��9bHR�����^τ�
֊=�6i���J�x�o�M^m�$�ԣK��8:���H饏��=B,��zz�5�
�\AK��!��	�\C¹��ʲ�)9J��a��5�ҕē�RhF��0$��|q�?��\�g	<մ�e�"��ͣ���[c-��^jt��$�)O�~�P���t�g Ka��={d[��|��^�eM \�]]�����*��/y����ݫ$�H�/ڮ��yA�	V r~�jd?w�K��~b߁H������a��&��+���;ޞ>p��3i�	���}��
�.d��J�-Z4u��% �Mr���ըQFV��'
��M����ɈG��@�vO&��{�bZ�Ã�0��^9�e����e'~����|���}��o��r��l� 6�S�?�1`��O��[��¥zD��x���9k� ��F���m,X`�/GgHJ?��U��4n�(�gy����� Q�hA���b��DDF�{`|'5�kLn����/���N��-���v��f��tS���_��r�C0~������ =���v7�Z����̏|�^4n/�@��G���>�1�%0��8�&��B���:����fDkcY�]z��I׀F�D��6,�-���4�8V	�vg�-����W�^巃�+�ཷd1|D��z:�Ne�\?��s�U��w��r�}[�-�K�8����/Y�@�aA�a�05v���
��~�����]��p�G/����:eX�A�k`�<ć�
�Q����2��T���)���~�0�n�uEwg%�П� Qn^�N�r����<����O��o�	���@�L���i�a��?E�����O��#bH�P�\����@��Y�؎���������1��Xw;�)��\�d=����7�P�S//�������׿�Dc�y�`~"��;��l����b�v_(jݩj��N;���^C������P�z�x ��ٶQ�V�A�E]�
�N^ّ�՝��>�=[���OV�?����*IՓ~�￠�j�dҽ����.,���X�):�Qe���Θ�Kt{�L=��9�G�p�r�~V&�4��Ͻ��&�����m �&����(�\KT2Z�o�ٴN��mɈ�˘c��z1��=�ɚZ�醅w��tK��iB@y�H'i�)�bI����S��X�U=6Mv1�>L  |�G�����e��B�N�V2��A�wE̺Wf�h�߾��CS��·xbv������T�>�1ne����N�,|B��~�\{��5�^���6P�@{��Zs�5ˠ[Oя/م�HiJHGΠZ���"E����^
�E��.��'�2Q����)�e&�mO�D��çR65�r��\��umF�������#��&�-�u�	�����T�kH/�<3��1�p2�O�v6�ݨ�q�t�uxHM��((�99I�������IK��:L�̝������-/�3�	��aE47^��_�����_���E�T[1���	�����T.!����[6^bu��
Vw�4Eg5�wc�[��g�JZȗ�)��F,�����@#�t�/o��T�+|g=�%r��oo�f�n��L[�)�.]�=k~q���1E���6�k]6��|�}"��ގ�'jj���I-�M8������-k�D �~u�� 1�x���e����PN��᳋�d�"��f� �ZI�� n�^W�A�V<f��C���q�;���)l��F�fz �Y�nҲ\�.���?�A��G�D��$��.��@2���I�ȫ��y�����������^V�g-�������_�Mz&�o�F.���|�ҔK6�^"�?J`F||���� �4/���j)�[�܇�I룚ۆHt�^ �D����ִg���J�JY��7� -K�T�R>�2�Ř ���;x�Џ#9�E��p�O� ��c԰�5$} �+���G�ި���ۡb'1�j7'��OQ.W�R>����\<���E||u�ˢ��K f��7R�:;�J�U��0�19V�� (o���>��'�\!��Ŀ�j��2$����ҩ���0�9CjTi��Y�F�M�*BӀއ%�*���@s\�WqZ��y���P� ����R��_���]��a�ƅ}8AV������H����u��t�]��Lu~���M@��-����{Ŧ'�E�̾R���B�V���r��CjY�Z������?��n�����$qh
-2"n�JIY�kWWz��_D��3��1#oL�i���>��eP`j3:x: �r�W�Go�xLKdlӡ 
�T�>��K!�@* i҃{�RZ	��l�<�+�uF���w���K�A�әS�"�?͟�&��*9�Ѽ�-acE���*P�[ Ξ6��K��5!�o�^D��ꃁ���;�^�ǑP*Yf�m���v}w㇪����FC�R,C�V�V{2���}�GF�:��t�q>TAʢ뀍_�;�r�n �沭�18)�5��u^a�6�ß� ˿�~�U4�IRx�.ք�VיEN����?
�����R���Ɗ~k�[rQ`��P���f����Y�Cj�,,8>�>�G��u�
���vEВo�|Ua���k;f$���jCӀ�~�����9����c�mhs���m%��E� :���/�N�G����A�(l� z�w{��+��?�_@}	6`�:��4A�ʔ��x+=hv��+2d؉рϙ�;ۇ�Kb0��f�}@Bi�CV�2�T����\q�Z�������^g`2+�(}���X�d~DV쇛4�a��B=W�Jm.�?�x��wOd?�!+첰,y:�#X1pec�E���e��C.��l�(��Q\*���+ܕ���&z�}�<G����q�� ��\�O�3*�Z�Æ��XGơ��ky�M�
�T��cmp�z�6��7�p�?S�J��hu�.��NFP@gm�����-*1�'�����i~۶̤�S3��97k���z��8!�Y�s�m�A�g��<� ��������Tخ[`�5'��},.��H®�=-j�|�K0ަ.�		�ږȴ���~�Zk=d�Z�fuA*���x�[����v(�/n��<(�%ԏ�ՑǐU�J<��-�"����q�W(�k��̖/$K�in�I��9_��US�f
��Y[�j�v�@uL� ^�(
�u&�� >�Cz�yIv,%
�l��IAm�˪�M�]�x¯��Ε�w�=�X`ҜԠYf���ɼ���ݐfi2�٘K�[xR�G��hb��@3&����h�-���pjh��ao{��XL�#wB}�f^�u�����@_����L�@�2�D+�f��8��L�&y�+��%�m�2�d���ԏ�{7�o`����E�=[E�?��9��{8��m�fA��;<<�2��]R4�� �?�Y�C�?�v��^�hj�h��z���[7�N�d� ���r\_�,VpN��w�S�Qb[F7R�Ȫ�����T���!��c���Y�{4YT��g��V��������g�˒��CUi�{���(����Zf���"'o"�:���0��̃d��b��?3��{��GÏ۰�T,��
a��eNp3D2tM�L��ӌ7b�nr^ �+����z��%qˢ�v��o�"��s����x�C l�K<۫Ox��z"�}J�8�B'Uܡ�4���)k	�|�2B�8|��������zW��j �8�߃ܜ�e�1��00�۩�7N)�U�i*� шO5o�M�Ձ#���4�a?�����+�u&�ϕ�	%�T^����d5��Fa���}	=z\�l3dvq8i�S�lk�U��3�S�k+x7l�/��ɄEu,���h�m�3�b-��:Rn(���D�]%Gd$���m_k��H��%�� �GN��v��&�G����Ϙ���k�4��]�힏�A�c�}�h倪��s��&(���A�"��e_�ǣ����N�~]P`��`qș��3n�������Cg��c�/9�GY�ͼ>;�����< ��8�+_�dpx��Y����Lp,�a*�)�yv�.���!�"���U��D?��y�cBë���$t^���h���<����8�~������ջ_�.�k���+j'�ex\E�~ܢ�Z!g2m?�Ǔ��f�3T�ɋ�;?���',��=]��[�P�X��ew�)��+��W�S�-Tv8���ٕ=��Q4�0�[�a�q�;P�"�.:�~a���K�M3�WZx��d���Yʬ�O�E��0~�YU4���By�8����lG�n.�^����K1sDRJ���/^,�{���~:8Ea
�IkmxK$LH\]g��Aa�,R<s�ku8����U�[�1.�y��\�'����C�]?��3c	���Ac����=���F���K��j�&~^R�a� ������ �w{�}	�I��1��l��z�s���a�c��\DIvV�˽ů�*�xkWʪ�y�����Y8'���b��s�|����mUf?#�Pʤ}-�����'�c�(��2�[H�m�U��|(���y�����-)� �+�2{:�1�`�V�E�$ ��7-�y^������&=t������ecn�Q��D������L�������;�iU�[o�&E���?��[[f��ߚ6�Ll�4�b��,�b���1B�f�/�.9O���b��J�2�<a{L$t��)�ㆆ6�w�.��{��b��h�P2�DZz�j�\�?5$Х+~�Ŀq2z;��s�ҽ�P;����u�h}x���a�Y�,Lp���
 �o+9@]\����ČesȖ��D�[���?��SdݞӋ�DM+�t��Z>��lC �!�qW��
���5���7�%L��N����>H{�}1�Ϙ�,	fɞ���\�?��Š��{A�k� �OPKy��Qѹ�rG!��TC/\K;u��ŜЀl%�$��K�#��E�
��]�M8��\���Gu���7���b:O���;w���1��<��#��%;�G4Y(?��LW����J�l�C�E��X��L����Ì�����b�������R)�M#�=���,��H����*G�F�.f�e�z(/�9�c� �a�G�[IX_a�=�@��+�F,A�)s�W�Z��r7�|�W�[�K��ASq(d��Wm7ٙ&�Aps� 줶�	��Oy����1��,�E�E�FÞ�~^;c�]��-����
��χ'GГ�.�@Fs���d�r�@��8��Qbnyj���yߙŨk�_;)w�	鸴�վ��ih�4.j�@��Vw�����=`�C�)�(��/�����xH7��P0Fq�^����b���g&l~���tMrY!\%��Rx)���y�)��u��i/�evʠ�-�;��6[��_S�5(��m^��HSW�\!~4�-�\��=��l�g� ^7��G��i!�B�H��$�h�4��5��+��i9Ka�޶ʦOz~�9�`��|��3$��^'�iD��,H���P0hT�i0�����6�iqH`�	;�w��yMI�dDK�_e�x�2���=H����2�r��*��wL�,��6HX+�m��U�!x~_uR��U'u�ZN�~A��N|c]�{͊lu�DI�^�:i�Q���͇������U��~��b.wuw`kc�s?�uU�$�����S�b���a��c�ڲ �<`P<��^?զX$�+���)md���2$j�R(Ug�N>� *��(��o�0=͖����WYwx�I��b��x=Z�_�bK�i�6 �?�I_�.�\����D���j���7ؗQ������[}RE)�����cB�Z��t��ߴ�i�~,c*�پ�e�Jҍ�1�Öw~��Z�eO���ͦ�^!8�W�����>7x}��Et�t�s�۔�Q+��?�K�� �"��F��4�SSf�T �'M��)��=�c�h�����E�9֌d�*�Jh]�k�� </��{�#���j�zX����y�����N&��<?�ܯKV~A�1��G/4�y��TJ(�7x�R��V�w�)V���+���}֧�]������E{�ڙ,ꂔ���׌:���4z��zS{�^��y�J6���=}���B�����^8AH{#mb d69�,"j
��"}�ﱖ�J	�W��x�`f��� �UF�?�8��ө�'��Y��k&�ҖvoЮ/:�nŒl�u���k��[� �d�g����[���:������gxa�׃�i�J�������IG X�߇� /��I��G,���C�ޥW����O�^������25\騈|�Ŷ$=F���9��.�j���@%l����Z�VҔL�cW��Ƣ�w8�h�����g,��Di���.Џ����Hb蛩&�r�{I�%ʭ�~?�@t��*q���lN���Fr�g+ ������Ec?ٴ�#f<��3���(&�%V����"�����
�{"-�A!ͦ���Po�"x)���	I�Yg+���u;����8:��G����&iT�2�}�蝖s�Z�|$�u�C��Ty_���LM�O�>3�3(y��{�O6X�\s$i�JDgr`��Ѥiq�K�Ĥ%�_��j:��oc[�&v>��b˝'��Rr���uE�~�b����@LV��J�5��}�U�b��N�an0�<&-_\��gh����g���&�U���C�Z�#����tl�P�"	�m�9�V�����[��v����~��0�{�� ����H*����W���[a �ZQi����,��{��B^_|8uF��=}�pzB��)~�M,�|� ��q�ik�}�mL:tb����������e����}�0��,`����)S���3b���x���	�� �.���\a*�6
�8�M�FN��� 2�׮r�;~P�D5e��Y��#I�V�~2�Պ����i������ޒ!�:9�I�����גB�����9�GC%�θ|�@��5�>fu?J�Fj+��T�ؗ�A��K��s���췐ЕߦQ!��������y^#� ��h�K@vT�c��,i�3UyPub��������;�#�O҅z� ��ͮB��t�)���#cˤ���)Wg���LL������3G�$���׶*���>
˛YɁ��:ޡI� u��1�\ylA)����F�ƌs%N�-��=��P��>a��q�ĭgF8������y�↤~-|��E]yơ��.y���sl�Q��� ����-�6T$�QE�966#��=5���e����;
H{���TY��aƼ?�b������"���߬]�@��{��a	�q\q�e���É�YJ���A��(�����6g].v^���j�����~�����A����C��nQ��s��������놲i��k�^|�P�T�bǕ(�O� n:� H�Dz�؞��}ʘ]�pID�+��":o���KoI6����@_�^ZY��-�"/U�\ްeD�_0N���'�H�*�T�nji��w3Wj7u̅[Y�ӣ������me�bJ�Q ��9��苜
�?јZ�s���	��R��o��[َʉ�s��N�!��4g��O�i�z�Hm���7DM������@Z�N�n��U����e��0d����'F����JKK��irgk[)O�.kT����f�D�+nM�[����r�^��V�<�����|8���U�[��mj-�U�(*ȷ�*'Ɔ�T\1w�겪�-�6� �.O�=���� ܽ[z׆�����H]z�+��G%��8�#��ە3落�`D�B���r�q���+y��dAQ���!���
e��;�Kw7�(*�m� M]��-�3��ٝ�Zz}m�����;`�O+X�2a��P= ��ϐ=�`����.���ڊ]��؜p�����ߥ��uH���Y���A^9c�[%N��5�>���'��K�Q.�����^V���������N�"^}7y_Nw��c��=��f�!��Ɍ$����|�����?�C��g���5�0�.VNKe���B7��&��������ב�?:�
lE�z�~�T3��b��E��jn ����`�H�2��{A�U��i��		���V��Rr#>��W�fj
�3"z�X�^�s���2��*�&��"ޣ|�6=M�.�����݀Rv��H�ѮQ�3.5^�NΩۑ���z�!�q��&H�M;�*{��D�HN����g�H�̝Mw�J�<��<Nu��r�|����0Ι���JBM&��6�p�G