��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���,���`�Q �����6�͍	),�6�md|_��n�x�"u������K �5owJh�E��qڑI9����%,%UEwf�x����;.�9��p3��,/�֤����"��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>:��cG���Up�Y^����˚;���"J��+��sc��Y6�f$6�5&���z���������`dcR�+��b\�v���D���ղ:h�W��j����='�5Cq����7�r!��:l�6�Fo���_˪��k��LH�]!��0�5�sֱ��'��!]ɻ���"	Ag�S�#kq���,���TN��#t��`|V�u�m4��0�c�WfC��� ���� `��ɂ��#2&Mpy���v"K�/KJ�ֽ�jw�Bz|l�#%�ȁ���ۻ�M1�t���a
M�?�a���t;T-kYޔ�z�[˵,�Y�Pow��P�+�_�2�.�z+z�A7�}C:�J���w.�_,q��xLNiP���
q�����R���V΃�n$Q���� L�'횸6,��c��lN����x׺��%��_d�����JQ�K�/�5��N#��Y_�Y9������ۺ!��iB����4}�0��a����7�����a>m�pJ#�`t��ąyz<m���� �O?o�_�έ:�	�`�����즪�Ϯ#(��-0{nb�?��{9د�D��#?8�O����0��aX��_D��p3Ǹf_��=�dԮY�,p�p�B����3"Vnb'7P��zT?��$d4���_ՕG"��GIT���Bꞓ.ʲ�������D[�{?����Ԓ�~D��)d̿�h�o7�!���sn�	�J{)���Z��v��߭��ّ6kf��;=B��;ᯠ-��ǻ4�v��|l��ݒx#��֑�[����U�~� T�0�b#�E��I�*��Xd�
���t���
���%[���ҿCNQ�i4J�`��C�;��gػ#LFt.u.�+�\�HM��cЎ/t��Q_~��1�I.;r���;�	Ǿ�(n�\³��iY���2~����)L�˂']2�H.&OE������a�Ȑ�8�4�PC9uMP$*R߷�8t_`�m�3�C̈́�k�w����-ԓY�n�qu-<.����V��D�MV;��'Q�f�	�h�=Ub�_@�=�T�H�JQ��5�|������U�$)6�\�̼x|!��Z�O@n��+����
H�+A�-$[��ğ-���h���.�O�=�[���Y�P����z���	�c��ˎ`s8:.�C�Ń�؅p	��"չ]�<g�Rm�F�W't��$IFkD���3y�32	�X�4����&���srܨ�PT�ʞ�袼O����	0���K�蚍d̜KZ�~�c��:���U�8F�sh�ܦq�#	��6����5��j��}�X��9�Шmv���b�$��NKX�m �$v���y�炝�7�����e��jRJ� �c��\��@l�4�s���jZ��"4Z[��}"�Q�5�P�*^�Ų	��J�$�J�h>o�o�\ ��d/.�,������t��IOVI�OYfK���N�\}�/r�I�O���ʇ49^����%������N��������n��4,����K��� ���d\I������7a\)�C>ȕ<\�w!uF��SOP9���.p���P��pemm�V�+j�1��%�b���:UIo]M(̙l!��QrމS�=����G*��&wr���U(}x��l|<x��%-�e���%\�*T{<�J�N�!�2v�t��>I+�II
S�x��^���SJ#H��/�6G���WB(=oTi��!�ޅn���t�+�T	֒��B��v��OG�����GT_���|}�jC�3��vB5�U�jM���b7��\R��YDEa��\iZ܎$J���(�7�X���4=�a�&��(����n x�0��n�մ{z�E�٭st��EqUȻK��H4�AƭJ�r>�qUۓu
�-W�'��|q2Y@�����U8y�<���;zڧ<d��;,���"-��C�u�\7��e�*����]�ݩ*n(�CL�3DG�r>���ɵ��/�����U�L��)��Ж��u���d���/���.ckl%8�]�����_����=�v&�.O�.�$��l%i^ڍxQQ�dc�
���&B(�zS����N��R:�5gd�ءYLD�iő�ҧ�,�{\�\���E�HeЌ��5�
�+�1��bc�2:Z]��7$�0b�P�i���@F�t�)ݩQ�vi����|
9e�G�̆��9�2���A�p~\�\�c��\H��^�1��^�!���)�Y|	�jr�|�~'�����jdh9�'����&�|}��[�f,�Cɭj��m��v��� E(-�w���C�JD��G��X��
�B^p�Ω^��!�d攽������M�;�����S�Yc!\���+��C̬�=��Z��7�v㭄�wݓ�۸�E�%��C�,���IEo`�]4iN��>��)�E��>���+�.�zФNCg든�H��{���S�����|z��eE�W�8��@=1�"3�o�BʊN:�6����-,b���9Ω��cU����Y،[ ��:�Ta��6(�&sW�/��SO�p�$O𒼊Y��vbC� Ȧ��(�4��T��᪭+��)���2�"� Z9Z��إ�߅-���5ʹ�r|4���=Q2	�)B���bI��Յ7��,!]CuC����I�nnW�1��tK�b&(N}CC'6^��7?VLk0	`���t��bci�����*�p�	�c�4�/�u�SQ�;�&ʜ��������I�>(�	)'���5t�7Ǆȝ��6�|$����pQ�У�l���c"��<��9HU��0���&N��(a��cd������xŖ�@��:s��;ϵ��O��[�5�r�
Rwh�gQ��$� ����^�����q�r�|�D�����6�Ϊ8���:�{U��-��:`����K�b
e1u	�$�D0-�n:ŇChu�m�5�ͪoluU�'Z
ԑ>7�̽S���;��E�K8��k�+��z�`�d� �dT�ʟ���w���T�]�m�l�?�ʾr5��w�����.5�i�ȱ�?@�' �Ã�9h�I+�â	�(M�V��VWu�_x^st=go�)���wM5g�稬���r/��������v��1��p����A���W���@V�?RΓ�E	�o5j��3��tpo�f���ս�	�2��0�����s�L���"JLЎx�F��8����ƀ����x��F�I�F���Ѫ�&T0��A	���Ɏ�=	�Z��*�@��0Ϛ�?L�їq���O�y�%����%KW����G�Æ-QU��y�)*Ċ�w�r6¿yo��6R������6�Yj�JO+6�Iţ��D}�)m��Kw��ۨ ���eH*�c��_f0��W�p�w�
9��_��P���6��=���9����W����st_Vʓ�x�{x>Ҳ(��F��ME�HỌ�~F�K=R��׆PH���tHa���K>��"}�zB�]^z,Y�nn��lf)�T��(W��^����X��1+�1�|>�9F[�Fb�f������v�9o�#K�Y�j�:����� Z+�^C�>e�(��
`�5a�o��6�B�Q��$�c���������g�jj���]���z��X{m�6�R���8H����#�a�pO��(��B\�F��1�C����M3�VU�7Y)ҏ��l��cQ�[nq�qFT����O(�ˑ��=7���m���d�dSŠ����k�T"���<�G�x�L�t��:�gO����E��W��ʄc�ԃ���*�oG�n�Ѻ�AR��f�q�T�<@��*j���Q�SE���{�V��t�>��C�)��?��^JФPek1�b9r>��?g�~a[��v�;N��^-���q�.fK�IWe��� A�*�zJ���LZ-{u�yƨ�ͱ�T
_��x.o���PZ]f+V,xxm�GɹҒ� �^�-�p!�a k��gR���Ym]�OLH��p����I`X�ǳm����&��[�@�<osF:���`�yl�E'�@���X�JfT�{f:�d^F��}D���ن��j?eh�^�϶]5'��}�p���I��E$J �M�Eg3 ��ⷎpb��e�[�4�ܾ��7=��0|%�R��cy��(�J=�t��S���F�ش7X��,�����4��U����$C������uU!֗=��~���g�:*���X^�{�Ć�g��gl�Zн-7���1������5��OU���f�|�ǫ�zC�	��ՋEJ�r8Ҭ%����ᵏ��aJ+F���#?O�v�}�G�.����\'�:��jR�#�*g��6����N��L3�q��#�e��:!9u�,՞�W��.���Z8�J�/|��笻B�6(���]��(T��Z����֤yԆ��L�qJ,��&g�J�=Ԡ�:�Z�:�$f->�f>��3�i\�ۊ��9���,6>��pz�'�Iz̈�(���)	@����G����r��$�ݥ����]��ppb��I��۹6�-��j:A�L���y�Pqc�E�`ɭ�?�J��]-�zx�b��b�SY��ʊ�W���/q= `W�_(���-H�GՓ@(�Gٛ���Q��k�ֺ��Z�8�(t&	���!8��6Qh��ehϭ|=C HV��I5�9D��F�@����D�{9�֍����uQ
q��t�t��6�����&{q�����HM�\`ئ��}��飶ɌQm ]�k����)�o��hAŶ֎(&����?�\K9�\`~�y	����y5��R�e�\j�Qo��*2�q+�\�0W)at�G��ߓ��lZrό�d2����\.�V�ŧ�K�0������R}ԯ��^�w�e����� x��0�J^')i������@(~�?%�ŵ�P-��P2��q��҅ft[7��PPuW_HB����K����9�W/���5fӥ�IC9v�� v��)og�����\���ŏ:`D+�t-�	�˓�����oy%4;t��MH��oa$�������I�u�Y]X\_ ϐ/�d�z?��� ]���v����wu��F�_Kz����Oa?�sb߇>b�ڕQ�/�٧�ډ�2��TN Y�w���kU��O].n�������5`
�EE�!Iqn��xUj|W�tA���s:^W�i'�[��S��ױ�~��t��ˉ$o-� Z���)�2�	�E��NѶݨ���@�dQ����H�3q��}��U;�/���j_�ZZc�.�;ł!�b�6P���jP>]�=9���G�O�k]0ϵ����T>_CC�����O���E�?����]�vOS~}R9�@,V~�"d�o�g��M�Z����{�q���ڝ/�j�)"���S6w'3ܟ������ C#����y|�fڋ���.N=s-3JUT��>�eɵ��)^������ �ô�Ū�l>|.z�ȁRB�I<3X�lL���%aX=L�N��6�A�F��A{���{KG?�����M��_A�pm��O��&g�7�n��mmS����%/�)�Q�"��߄���:�M�&g�ȣ�LF�S�vC�ߊ����� ��s�GT�I@����k�smA�D)É��u���i�݌{h�����{�6�-����f)_	=a]<��H/�{)�lA)����8~9�/P����tf�+�������������wǼ��)TJX�o2����5{kGg�o��N�<sf�7\��?z�~�3�Ġ�J9������a�̊茳)cB�g���LYb�H��NN}��4<���Z����K%��۞L�>5 �vzh+~�視V��|�.\�:�O�U�����(��a�᠙қ'��������h>���?ކ��xJ�=V�P���I��Y��{z�Ԧ�N"��:�J=At�"y���\6���.���~3����mZ�ah���.H�-��$\������KG���©����/�-G{a���S2லq�� ;_3@ �V̗���fy��T��{��8C���r ]AKD�c����~Q���q�`����H}�G��n�O�VD<#7=��;��˜�5r;�/e�����$j=�	ȸ:J�3أ��f渺\5U#�X��z�s	�a��8`X��	e>�����@c�uKWv�� o=�N=��\G����$a��V��mH{ (d ��BJ���E��7���PЬ+U+j�"���"�HhgǗ�J�IM��$�_I	������:o�l���N5��v��c�	�(�gx`���la��������+$�:�<�>�iKv[h
"���ңw�5W��n��Q���!��`�mhL��l���
�iCK\�]�e�fg���t^�c�BG��}7�Kkf��~ox�f+�(ƈ�1D��t/0