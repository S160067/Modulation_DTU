��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����0� ����遼�6������"���#�{A���'j�Qj} �}xT	g��F����a��f��洜K%g==�Z���L1������bG����XB�k6T��w+F��3r1#�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>:��cG���Up�Y^����˚;���"J��+��sc��Y6�f$6�5&���z���������`dcR�+��b\�v���D���ղ:h�W��j����='�5Cq����7�r!��:l�6�Fo���_˪��k��LH�]!��0��-����{��¯d�Ҕ�5.��s�ǒF�C(L�G{�Z�F�%�x.�M���L���³�Ą"&�5"���Z���Ku�@���.?�DL.<��ײ����� �vW���[ ����N��)�"��rFc�B�F#�������~���
u���7ǉ�;�o����ʹvCZ���o`Ä��rg���5/f�+M�y�ؐ�?16)k�� ������$���.��MԞ]ekW��%}�QS�#vm	���0�3ժ���;���0�CK��{�J�����v�h"KX`M(;I��(�az�7:_�����/ͰV��t���S��<������![g3/��0��Jy?{\��Z��`O��-��',������K�*>i��Pb�X-�7"�#�$���ތ�4FY�5^Nǖ�W!0�#����`�h�� ����x�V�Mc� �M8�)��;xS�Qb.Hıxt�)��=����y{���`�4%+f��&]9�����RN�7u45�v�}@�3�Ѩn˞� ���R(��SO�i,[��%��݆�����p*�f�����
���ʺh[�i����i���� W-�dW!|Ũ�DJ�hF�JV]��sv&�ݔ1ƙ=��a �j�0f�a���c�4|���[<���}p���i�\VC/{uRS�]wV�<$��G�O��j#`�lW���=V&u����-��)����c��mHR�O��3�6��2� 8'/��cŐ ���O��:�FC�C`��[�ʶ��tp�:�1�Y�@��G��b�ܱO��\�/�\����&�5S6<-qU��O<Y�Myl:O����b�sv\qr�&,ru�`�c���#����G�6=6��z���P�19�]�[��<`WwEHص�,��������.���2��fq!*,�{)E��	���K�S�Ga�o�o�!�W[�����3��>�ٲ����Ҷ��sk�����stڛY�NG�8}�!#��5��;��1����O��*�l1\�K��5�X9�@6�![EE΁٫U�^�-�co����X7�7KCwhg��-��O��3��G�7]��5C�L�0g# ��w�D$��	�7,��xˠ��~X��_JW�l%�V)sW�s(e����~��r'�&9�O���P�U���p�|�<����2+�3%�3��Y�ydC�� 5�"&��ܲ�|%�]x<���Ǧ�@Lq�aP0q��"��n�p0���,�P��q����)W�["�?��y�/���'G�ְ �L��+���F�N	���rl+-�h],V������	��qq�VSKo����>��<��� RH�א[�|��&�������ͥ��P�,�F8�e��ʺ�/˝ N�f-b~s͏S�h4��DנGe���e��>����^���^������i��@��<���HګD�{~$�Is�Xm4k��L����m!�@dBO�sZ-K]���~��vm0=���܀��Nz�g���!X��F�۷h�5�����
-c|�j'F��Cͧ]we苂C&54:,�T��=�a`�Z����fs���`��ɏF��;��I����������,�o�����HV��a
kLР�C���i���ͧD?������>'TD���3����M�#c��9���3�� %Y� �H>�=>�Z/��o���!�ɭ�k�=���=��S{���l��z�a�{21|z�VvE�tM���9G�#�c�� ?��B����O���bQ(���swv�2�ϕ�$�.M���F�^f�(�
�L�il����,>������,�����j�M��S�r�>�u�O��R�P�P�Y��:p�55|��WQD���8��z.�Qt�h-�h����#޽i>)��+�J��'OXH=-r�=f������x�̭�(�E:�]��U)>��G]�M$�7�M�;������h�h����f�B��r-P�*Yq�g�߱"6D�k���<x_���!��7XY���:�$����I�c���U��WƼT�i�bAo4�hXY���e��DÉ(a=d������{�[u%:9�������M�}�fE4�����װ��*�`W�n���kB���l"����Zʯ�q�_�k�Χ�����05���'&��?��D���	R�����#l0�t���j^�l����c�R��a�T�`>-��mէ)��u��Z�Yވ���|���uyK�D9��*�:s�_?�o�g��ٙXe��W���΄�ЫN��_p�|�'M!/K�e.����MS�v���#��s{h~��r�}9�4�-'�C�x���]��)N,ϹB4v��{0m�����VX ���{���m��{Y\.Ea��N6��,����a��Ź`p��N����b�v�����������B#����-#P��E���܅ՔBWv����*�˴�M�N�!.��:�?���,CK=m�`�f\��C�~O��߻K/����b ��J=��� ���ʕʑ����dT�Y��'�
JRi��q<�4�� m֕�r���~�D���_����)�0{��h)O~�����QB-���{�Ì	}F44�	�N�	/j$$�u��>�dH#����4O��C�~?z�lw��X��ɕk��^O�v.TC�l����]��@l9"	w���S
��ec(]w����j����L�SZ���\ai?8DZp��l����k�М��7�z
���`}�0��9n�rsP���9�m�V8�Wϝw�����4r\���_�N�`��sҼlf��`��3|i����W�p�[О��.�O���nj���������d����d�28�N���ח2�����6�!�� �k���N�|���p�Pz:�U��S��^T�e�q@LH~5\�{_�4_���X����.��g�W(���af�{a�O����F�� �0�����-G�-MH��rH��ު�� ��:��4Ha�A��_b�`����d�����~u8�X�u�"�u��A��X4�	 �mҥU{�]S��l6S"�j�zM�CDA��X�����������izf԰ �U0�M�
|S�^M�&id�.z�ư�JPa�I7�v���X'_2��?.�o��@�n>�<�zB~���6�<�G���T�MF�@r��E�:���yI�(�O�Aj�jA6EE�q���#ᎂB��Q"���le��Y�Q���p�̧���^s_y�T�[�т>Y�xI�N$(��1�.[�I�[wG�$p�����p�O]������y��w(��d(��.k�, H�`	]���S��=�e�R��B��qB3��S+�Ml����
 ������|���y'�4q���k?�X��v�{�	�P�s裞���z�S1�o
���_�z�D$@ˀߘj]	�c��:�i*�O~�tMQQ6"��wC�uW��m$�r��i9��Qy �|P�����Tc�9�$��w���|��2���/��a"XA�5`ǎ�:�[Ұɇ��BFZ����d�/�k'��ʙ���lb����$�
$�Gg��P�G�ȄP�aw�����c�>�8
�x����)��f��C�uO��v~�pSv�}������"J���=4Z-��Q�Ra��aqZ"I(�{���D�y�^��K��X'W�h[A����'Wǣ3ޭ��[��vo2a�l���W�*;�� ���L�_Ir�]�GǶ�}00$��*9{p�\S�F{-�هo\��,"�G���?�?��:A�@�{�(��5gDΐ�H��.{�"��D͙���C�rB�U>w�1n��a�g0�z `"��¦UTu1�H�+KA&vW��Q��o��<��[5��?�8����zK���H�\Ef���^F�cAO�HV��`Jϥd;2 wx�2�+�5�֯4&�����t�����+u|f�D�����FNne�0�A#�ZR���� w�Z�A$�Һ4�Ġ�rVD$���0$S�$4K��1�q$���V_۰�{{�7X����c���G-�'�:R>r��U:���"���e�BY� ���X^�0��N��� Lj�p�[�`�7�����a
���\��D�4�_3�*�z	�wJ��4��1�xnp�*	J7@Ң�i?yW	G�MI׷z�>h��	�I�I�v�u2�̹i�CߨŹkt��f�_��z��߷o�ص�<�8�\2a~�Z'��W��Z����D�� ��ØlE�+Z��N�\ܯ{��nh>�SCg%Tf���Q�S�L���0b�	ډs�(ܐ&I��;���1����is{�b!�$����H�{�V����'�)���p�&LE�T�������=����k�Z�֋J�\��<�6XY�������o;��#o٥��8��`�h4��������5/�iA���_��ԉ'K��e����[T��Cۨ��OZ��	�����(�Ԁ�h���z��t��n��n�cԆ�F�xƻ;|z&�^��h���$F��r��6��%�d�^/ V�{#>�q8�E��E#�8��+N�"$+��qG���#8�w�aT� {�� ����R���t�+S]� n�p�n��*d:��A]pLρמm٨��3���g3SuFK� 4�i�b�N��k,������\�z�t:��p�����7�kg4��Z ���7��]�mc��٬!�-5@�v��`���&���c���r�W[h�R\�
���Oq��i�T
_�0���r�>�L�}�њ�ƌ��oaT�т��;�/���J �j��,f��Yh �5@X"�]���q���=/)���}�O�н���)���pgt��/�4�5d�G�����|6<�Km�&%��ГFa�v��K��)Ѳ��"R�S[΍��j����I�ɑ9sm��'Wm?۾`�F����M5X�%`��⋨�%Bs^Tn��>�VR>�{W�	����;b.,x[\�m&�q +r3믭�������G��R­4BV�'aR���B�	c�i�x��85RSL*��+�
t���s���+����8%��ϔM���.�؇�&�/|iy�X��h~R��ǁ����}�Jn�x4F�g#_��޵X6.�����w����/�&]��K�	G�@�4rT��ӵ��˕�t4�`Ju�-�<"x�0Oiǅk�� 7�NsQ{��н�1/W�!��,����3>[��t]0hl�NǀR��D�q�����m���ﮆ�[����4�1cE������w��,#�]"eW[X�"�OQ� ����s[`�.���4���iG���g� ��}�4w��k�aY�Ip�ה_�jY�V'w;
�Ѵ(l��4�(��p�n.�c3Z����?�����T����F�i]�?������%�2��V�%z���VʯLTv�NJ9��#�"�w^���c�GPx��X��c|�Ju� ����B���i��SJ���+�'����V���9'TM����J�Z΃��>Q����@M(Z8���&�Ο�88�
��M��J
�_����A! i9�m́�u\Ae�ק�h@�'��P���u�0��.�[�б.��h�y�z���T�*��i�N��[����2#ɭ<�~�8��⬕�i�pY�@�ŉ5;?|ѣ��ȅ �U��Ǜ4y�����S�w΂B�N�jEI��q+_��:��v��dK&��$(���J��p�I+b�?���"]������6��o%�ӫϴqOtῶ&An�"TR(����	�\m��,&EІ����S�˶�T~�7���2�/Yo�������jc��+ެzb��0"���8�6>/ݴ��� }E�?a.�k�2�D�Y�4(����An����$B�Y�wE>��p���R���a&�vdT�ݽ�"E��G2ST'
_�+���$�®O�i)ݔ�� M@��7�b�c%捦.��͸*�u�����k�Mc��[���Pc9 h&j�K섨�@4���7�1�q��ߩ(9���r�W��F��偿���o$Z9%�  ښ�U06�J҈�D��JG/��M:kT��60��=U�«�s:Y�ݫ�܌��)}�m3�g����}Lİ����]y�V��a�37vGiz�L���9�\=V&<#��|ʆ�p~}vP8��R�ުO�t�F�|�>M%���7���'׊�