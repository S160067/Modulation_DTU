��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����0� ����遼�6������"���#�{A���'j�Qj} �}xT	g��F����a��f��洜K%g==�Z���L1������bG����XB�k6T��w+F��3r1#�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf^��$�i�g�Wɐ�)
�Ql�Y�+6�iѰ�^���d�u�.�Ye�ZG�$*�f�pM��Y���f<���YB�H6]��^�8�G{��:RjeQ��2
�ƣː��5JLO%/.�)����\�
,��YIw_�aJ�/��]b<Q�	������*;�ե��O�T7�f롐O]�ETt�ҿ�aǥ�ހadz�)O�������U2�<+;<!����ֈ��}��,Q�:t��9�ɿܐa��c�.�Tp��I�/��ekS����V��K^	_�����q3�؇�Ѝ�Mx���3�6��3�*�O;Q�Ӊ��	����+&����/ƨ�KC�apd�a{�G>�vc��a��l8�i��������Mi���8��M]X`�Nx�c˨��}��Xp�@>1D_.�>�T7R5#I�u_A��H���'gel�S:��w�����f�s�7�~T��!�o<�-�+~'��^B���d������9���O�R��{�h��� ����FM^�^�d��,�S/��zGR)�t�G�PO�_����͹_`a;Z�8���|��$�d�/�AV��݌PI�?�,�m�_цa�Y���RG`�GX���zk��9���v��l���n����P����f����h�jW�^ ,�{�7T�e���]�t�x洂JL���o�KT50��L��a��P�T�Th���L�����@h�kR��V"�R�C����15��
�i��N�%P2<�;��P�:1����li�kB� .��L���8(;-!�����[R�1������[��l�v%�&�NFP��At��Yr���"{%ݺ<o|�W}����������_��t��\�sq�3f�"�9�K0��-�Ok�eN��D�|>Ĥ`Ɛ�U߬�@R��njV#v[�ن�%/}���f- ����8:��Sz�%S4���傯c��"�K�ÇV&����F��ʵ�'Q`�uQ|�)���ް=g)�~U!ϩ
�׫p���S���5ӫ�(��"���z��)o��²Ý�SR�g�B#�/J��ʨ�NVխ��h�PC�I���G+������]H�R���a���'&Ɖq��?G(�=����/�Tr�/�z
�ֺ:�3����*�J>?b�J�v!C�C3v��:�,;(�Q>%��tNX�#���|�l)�M� (���+���w���|����k�sҳ.�:�r���O�1��2^�J�IׅQ�(V��T ؜(��[zc�+�����}�z���ʜ!�R��\?K=X��#�621-{%PנT�F��ϊ��{��.��Ȉ[u�a"y��I�ߒѻAw���ԝ�q��NOYj�g"��թz�G���_jZ�]+����a�陵��4uPʷ�&E�k�r�l�E\9^�y���q���\�i�"M4>��ND2I9�Q�3V	�N�h���0L������f�u: �s��Y\��dெ2KW
�~]���s �%�����Ԑ۽�Ckl��|K�&��f��ܚ<8E���u�]�\s����1&L���gwo0
�A�{���9�n�2�cت���~���m�B�4oy�����aH�W~`�Ms��,��W�a�`��SZ�V��"��4g���㟄3`=�]�^�Zǔ�K�7\�{V��s>��.de�ՠ�XP�G�6H'ƅO�tȦFZ��A���fd���p�N���'������6kDI9Q�	J�+���j�!�e������O�>8�g�]f0]@ ��Q��c�C�~�5�7�o��F�!O��B��V��˔�γQ��Y�.�"�$:^��/�5H���P�_�%䜐+�J&6�nn��E9Ȕ����K;�t��+��{�:����A��<rv^��JjF�HBѵ�֭N�h���R�����{�&\��"��n��m��'��T�n�vw�r��{e	a����@���%�j�id@٪.Ԕȱ��NFe>,�����G�������.N����C�K��=m�/��/mH�ri���6�����ZW%�Ԗ�$"`��ۆ3JZJ2���l�Bj^(K�Ô��sSHM�D(q��'Nf���*�ܡ���>�_�N��(�U�j��hX�1��b��Z�"��5�P9���_5�#b��e(��t��^d~nhϫUkI_���5^в۱u=+\#;,7hř	�`%O��9`l|������'�y��3Q�ԥ�+���=kE��g	h�m�� 4c�^��g���$���/*��L$�I2���ƒ��dx7M�;!�襫Ɓk� �1Х��G�ޒ InS�Q�X9�=f��U�/88Ϩ,�����R0Ԯ����3��C�߸>.��w8?.oBf�'Ů)	9�D�ƻ��eM���gW�]�)���-�3�#��n����quK�NH8|_��	�ޠ�t��@3���>����Y3[)�%������ԥ�Uϐ�us��Xܜ�+�CzL��T���E]���(��z�r����X�z��N�OZ�2CM�%B*�Qx@��1> K�N����&z��M�����V�����$�F�l8�>⢴����O�hs�/�*�L�� �s2����{�d��Y{��/��A4�)��G"	�2�ؽ7����\�
9M�D!�r_�d�Ͳ���C��a��	�J��Q��B7 7�؇��������� fz�|��!�z>�EIN]��Z�؅�ff(ee��Z�R'�}��(1�a�7�&�NI�����+���?�k�=�
0+��H��B�#0�#�9r�����h�I���]��e��5߄�P��@�j$��X��&yUf�c��D�	b��$3���@�D靿��C1�����)3�Ω9
������2�i��Y��jZ������AukB� ��[�d��������z(2��w	�k�~ڠ��e��(/��ܯ��()��0�e��~��{�'��
@��=0���hMuVz@�Z�U��5㦉���@��&1�3�(�b�!v���_�ⱅ���x�����$B8p�qdS�[���_�<lir5fשZ�ʆ�����F'�	)������E6�ٿ׫6�w�ǥx�������?�qvB,/��2�_cl����KC�%\�1Z������P�&ܼ#��O����q�$�_��=+�<�
�I��!���_N�u��T��K9.	-��ۧ�p'~���<u�i�\����l�S�x�ޅ\Tҋ�`*&�LV��*S�B�V��P������s�j�>�����p��X�����,>�J�|.�<�n���R(q�?ƢgXym�����ކ�l�f2����5&È�TT�J�2(��C�%I9�H�u �<��]u�W�ge-�l9��򎂘��k�͝n�(]�
 Ǔq'�>i+O��6H�r��O�/�%���U_yc��<�5|J38�I��qkf_�cZ���@xy�8<mF�)���/+��D�$K����w+A��!�����{�?)��O�3G�5A<�qgZg��&Mwz?� ��8�����M���F�� �/�֧ά�6"��;�m�]�+�n�EQ��]O�Q�'��P�΅��W���TiFyJ�F3���RiL6�Ld��.Yv�m�ܺB���5�ن�!�p�%�a"���	�
�Ҡ`I���8�]'�o`،�M�$���ɨ�����^0�����FRã�x����3e<�5��M��v;{r�A�٣9��)/z�Ֆl+z�����:C��E,w�*�2���D��+�����营�jSүX��a�`�m˘č�/3��v�,��: g��d0�;ZBn���� 3�\���N��`�B�����1c��	��aρ��E�.&��T���aYuLߏ׎\e��r�}r��x\�ރҞ��\[�O����z;'��Ez��M��.�Y�K^�LS"��1{�89�Y����INu�5��f_�^�;��#�N�_��j�kf�3 �:�s̓�=r#�Z��s��l�b��b���lCqN71�\�������@��\�pH�Z��D�j4��U-�(�v.-���J8z�@�̰GI�I6�`=?i3dR*��BUX�C��h�������������|���Z.���#���(�=��كͺ|��&E����LM�d��u߽BP�'7��%!�,��<�\&�u�.>�����MU�v�KǞ�D�:�|~!���kNby����]5L����JH,�	b$��{���)��,.6~��Ђ����edB=[�U)�E�r"�c��*�!P�E���
nk�b�!S��E�ׁ~�zޕ� ��o�ߖ��^�pd<R�h]�,����CM[.�8�򝪩��� 4)����*O�ٺC�����@��������H���5����6�m���	݃���o+�>���� n�ʃ�C0mC��%��mM��ĵ*;��a�������Z�Y��`o��
�MJ� �d���J��uM�Q����./8_R7"-�!�)u�4��x���l��H�pE��I<;��(xw*�⋇A�a�����R0��Lέ���5�XO@�s%-���gkaC��-W,�j����`n��V�~G��N �n��m�_�������}Z:���D�]�JfQ����|o��S��r���Yb�w�G���|��n��ޔd�H����͑Y��S�\B�R^k�ڌP�$��$5�;s�߈����	��9����>�W������y�C���֥����Q��V/L�P��<v`�^�Qt��4z��e+U�d5�&�D�}�l0m(`�*���(��*&��y�g�]ǹ���q���t�hr����S	�񣞰,�����+�B�����Z�4��,C��8FK5e���^Lj�l�ڠ�������.�P��p%_֪�Gs�+�7H̵��^�~�`몫�DQ?�@��*P�?�ֱ����o���˥�ƯM�]dԨ��<&�S��[�{#������}���[�vYfSR��/���yG#.�D{yO�*�캱��bǘ��ޮ����V�W��4��K��?;K��[���x�������=��8X��q�!���?�W�P�G��Ma6�u&q�����:�"1���dn$U0��ʒBXv��a�M�b�yziL|���)��R�/M������7	l��#3~��.�Fs�#�.p�Q:M��b���1��+6�!�OKi��U9�p�e{|�|�=V`�'+C�ǐL,�a^���;4e)6�Z�̙G|��w��k4b�ڛ�!c-/�ը��j"Q�-������Y���%=X�g���^
�}�)I�2]Z]��Z����/��[��F}�^%fw��V�m/ۋ��f��+jc���E('�)�����Ky�/��7��p��:�H�P����r�㳬H�7T| �5F'cX���het�\+�"�f�_e5�i&<�~܍�rd͓n�|��B���C�K2���M|36�n"rx�ߎ�jC%6����ƃIg��:��HV	���?
)����aR$`HO2� 뻠v�K6����Ƶ0���߰�vd�Z����l |zÂ�w$��)|���L�va��$TN �a�����b JqR�c��fU����.�9�]���3��{��/h�˄Ow��=Q*x	����zﯓ5�Ҍk�U��&uS|�R;�X�Y��Lr�v��i�}��aKwlJXk�O�B-��v4sR�u�F��0�b�8��cRJp��]���4�_8�1w����H�����p�c�z�x<���+B�=����G�پZ8�rt���)��y�#S�-��Zm�Qa����OO�gE�W�&����j;a;�Zgi}�����q:��1z@0��V�roz$�-��F]����L�q��T��.�#�N�Dَ�R�4���<��&;�R����2e\g�?)?!�!�Er����ݖ�-�.+<�l��Ln2M���J��+���!.Ԥ���Du������@|R���CP�YH��L��'�	���d�ׯ�[jU�v�~?&~e���Ȕ"�&*��\B+� �0�?|n@�����b��@Qr;��
	��$��|�*�o�	�V�|�F#�'�����d��D�`4i�(�)�Xި�|}.�\ ��N�ň��Fț¶���wv�oKxR�;?5, �N��]*C��3(�m�Q���4ސ��`��tg�+F\hm(2=���J�_vC߂t��j��Q'��_��^n-ǫ�xź�#��#.[��T�[��PIT�(b����	N���(]��K�_T�\����=�����[Z�y�G�9<fBf5��!L�מcML�Pj��TR����w�����~ S���rTL�QK&[�(�I��Fr�!�S��sp�W]-;��������H��ȕ-���*K�@�|0���a��;�:�Jm|E;��|hR��Ji�@���>o�Gɽe4�z���M��%��_ɂ���؂^�;"~Qhv���Y�0�wۜ�&���|	~�3�1g���+�"C��qH[�U:��K�{�~�
�-�xI���Q�h����Vw�'UT��:�yc}<�Šu=O�7�Н�*s254h8R�*6��K�� �C�-��(��[��L�!��2�^���m#\�y��=�h�;�R���SɁ"H�~����lFt��z������l�-�7�b5����m���ԡM���(&��[WN��E���g93�>kS^���QO�`�����]>�jX�<Qn�"��8�_�;HZ�=�4#�����߮�y���uJc���<��B�\�Qn���~v��!U��	0R�Ԝ�� ҩ]n���L��@�a)�E?b�uws�
7�9�������1�y6c��m�af]��)�T;����I���f�� �&9(	w�h��+zz�{p��]���oL��n�z��6$!M;:$� �Ҡ.v;	�N ����A�w�d�r+ �H�,�x�ǒ���:��};��m���+�d�R[��
�Q�ƊN���V ��i�X)�p	���������8���ۭ��GS�Xa��gj�Eg�M���3"�5���6��]���2�Եdā�o�9��7V�5�87iIʵ1bS2B̬$5ד�$���1,���
Hh� ����tj��w���)�ϪC�v{���C��S�(B��vZ��z[�A�E �nV_��@x��O6�h�x�6	Y|Z�.���j���g]w��'�;��v$C�:Ȧ�eC�3���G�%7J��/#}H��)F�� ��]b>~WQ�����&��8��Ly��'8!>�@5���ݵ���&��4Uh9ϡ}�ߺ� f�F�F5]>���^�:���P\N���C8q/ |��.h��}RW�:�r�.>��u�k
�Z@P%a�~���u���r�\���$Rpb���ۋbAɝgS��*�k��R:��j�������6}�fT�"O�II�R�4��/���K��b�WD��3�c��M�y��n����v)S�-l�ʠN̍���`f��B[h�Ɣ��n<��u�o�Jd�]<��5󦆾��|6�%6,HQ?k�qr�g�X�6�;)�O!�GX�^�C��+�*�Y�Y��A�|^�=���	��9)'��<���c`�v9A�=m9F�"��)�^�q��6�&�3;l�3�/�n�����œ�������G������rpo���y`#����u(I�<�̏1]x@��ψz��^�c���)�����ؑ%��/��H�9�
\I�+s�{:Y���Gs�[)C~�Yy�Sd+��#	���.Tp|q�)�0�C�d�{�(#1�#�\�����7r[�Tp,��ص�,��Ϧ+ͺV�k<Tp)Q�P��G��q\����\눚ވn���a��g!%�#�X�����Hj��?c!,՛��ش�s��f@Җ��geȔ����$j֣��|{D鉉i���-ҽ�a?�a:�sNP��l���"�Xz���w=��g�w�ڡ��o�H�.a�P�.��i�����Dz�m��O�0O�bb[����i'��&](��f9�Ã�� /$ȃK�G���hG�����G�2��Q����ϱ��hL����"��ѓX�ԛ��Ujk��!���>��B7�$�<-�'M3�d��r�WBsD��$E��ЦHQ�|`޿��36���L(���׸̮���V���ņ	��(��1��z�=�CӘH1��6W�y�N��{A� �gsY �d#�,�����艐�ԕ�gT��2��j.@�4� 8����L{\��~Z1HY��C�</rV�\����̝�:��jt��5捗����nD�|7�Wb��zcv�����2i2�̾�z��w7g�nݽ,��6��4���#�ˡ���=V0���I��0ͱ6{�h	@@���+Ύ��j9� ��i31_�QQ_�@���E�;Ϯ�'<O�tc��0 D�܇�����ׄE��ź��!�L��-�g�D��Qd����YYx��{�)���Ic�#�]��_�̘�i�(z+'�T�1z����:E��mT9$<��[*�����?�M��3�=�H�hk�(��۰�C�p�8�P+�_X�4z��M'����Zl\$��.��hj<�4qe{�ME�vqU��y
�m�o��Vn��Һ�O��Pa��h�%��FaGV?`DC��P+��r6����C)pG�U��,�x��&3���z��o{��+\(LVR�0�q^��(�X�!�?Tt����l�b+1G�u���!ַ��ܿ�̸�w�|�ņ��wN���Jt)�@*a�@hBra�-Ё��s���aF�s��*N�Қbx���wSm�������"�EiY�z�ݖ�5�e��˶.%�b��B�h��>�F�(�����ML9���&���@;���)�b��W)o�N�q�X�Kܭ�YG�@��j��|t��,oB�Ҩ1=:��u�����rŘ���?�u?%愺�f���ZzZ�� �V��F(���ߎ쁛�Z�+Fv� /(��3�ȏx��y�l�q��.ۀr�t�)����쑁D��h�W��:�"_!Q$���5���x��</w�e`�'�����L0e���94��J�KX;��e7�VM2RG�	8V�TP�&����NN�V9�Xod���� �:�|LE�=SGީ$��=�K`�1%�_���x^]u�v�R#�Z$-jwV���T$'��-s����7,�4d�ã��1���*)UV\S0�̛����*g�h 2z��z�4b��)a �g7�ϵ%Z�g[���� 2��&�mUK�z�Lt��juA?u�vP,w	֝p�O7���̉�a��+�m���0��,=W�?u^��K	D�}���߽��g��;���U��9�؝�a��� �I�&�F�@���Ѕ{��t�#~��Vڽ���J���%ͪ�n*E8�	���z��.�;�!�>����C��+L�Z��{�?�p��v�öS?���~�Җ��+?��3��UU�D��!�t>�V��������U�5���[����E;��V3I��c�A�W���n��O�ঐk�'q��=�<	/oo����'rİF�G��o�ĕ��Nq,���I�>Q�������J,�@p*](+���	~iF�0k=�l�x�֑C���s!���E�GW�z`�0I�"���y(`i��ѥ�RH��p�e���|�)s���8�]��)�]/X�&��s�S�u5w��L�-AA�#r}�mU��6��]��x��I$m�ã\�&~	���>pv c�"o���ڴ�;bNF�C��T�T(���2������G�^Ƹ�iB
�#�z�����S���R��[�Y ���`r�{���e罺���k2�L�~�B_��(��k<�hf�X�Y�^�5��vM#.��Yl�!l_���XIl�]�J������B����`(w�Y����`��%����7��"}��&��J��f�3&�0ܜ�"RQq'��-�3�%.����w{?�A2�H:��*��+�����Y&ǵ9g ����,�~7/\��"Ȣܢ�kr��FUV�6�j�F�7��ʩM�s|H�#c_��h�P"Bk?�����,��zcp���U�*���a���d�F����zù��ՖQ��/w�ghCyOmz���}g�	#~y�'XjJN�������B�S���ޛ'�l�?�����소R{�ym��3_���o�-��*ŋ�`�%Ƹ�(�yްW]R��Z����a�=�Pc��R��m)s�K�m��a�R��ir���Z4Չ��w[I���W��[�2�b�t�u��ޯ;�-��	���)�ӂm���M�oE�-/�V�L��}؟�|�Ç�H��%>R��nZA��tC-DYY�uV_˿֣F��P�l�*F�n�[�>�"��� ��	�!�e�;�',�d�2���m>���@���E�d��u����s2fX�$R��5�$v�k�;��.� ��(�'5a���v�gI*&���q���J?�娫���J��+0�3�A�|�_;=��p|.�qL;!������T������#���Q��J���wU鮨%�\`%�Ŕ�E�6?��-��D=� t%s��ӱ�q�%���C{� ��[�z��L�Q`:��9W�ڂ08\�m�x��}+W>#��	��A�^����G'e�d���"m�Fo�T���5g��pE���N �Z]��['��+�e��\q�K\�PH#�<A�~֒�[���Ƃ��[	�i�a�q#��m���]��3y�-��5"�h�%F,3ꗓ�Q���9d��ϕ������D�	=^�g����RC���\<~#6T�2Ro�Z���!I�s�B8�U�i+�0���
��?f넇�3���L���/����R��*�����~d�b��|";2�4�}P�4�7��*-L���b˷U�'���-;�����9�l�b(�t�Yz�jn��2�p��*���~����uO׈ ��ٶ�,#�k�	a�N��`{U)�X���Q�,J+/`2·�p@t�Y��#��,Ty�u�E� ��?�*�Z~׸��Z���Ͱ�qJ�*�6|y��u��?�N/��J0��ƪB~���yt��Ft�i������^V�Ѱ��'��#�a��h�����o;�Ou�Y/O ���B> �~�|??��r9���oc+S��mam�L���Շ�{LrT�8���r�US��P@�^�*)��Rjj�;�7L��s�Q~��(�q�E�1����ZdU� -h*�@G]ԲCÔ�:�?�����_maO���}�؟�*ݗL����f�ۧ^�N53��7X��}'fPvc���e$�)�6&wM��h]�'�j����Y�
i����N��`�?�:P/��T��G�ؠ�z]ng�߂w����@�-���X������ �'v����8��Ac�K+_F>q(�{*�����&���7��\�*�^/nX�n�u�_�0m-��v�o��I�Z�]�wd[#��H!��1K6)�SG���܃˚rV�Z��K��
���=�L2�SqtEa�%����t!a��)	4Th����2"�}%�}_��r=�2�*�4*-�t�v�<�u���F��-��b���yː�*ay���M*��t@g�K�`�8�� �>�G+K�F~n��6u�x̮cbҿ�����@`8�f~��ɥ�{)���
KУ6��_�:w4��%`؃�����x��a�}�(5y)󦉑��"�u�Tm���Ǳ+�2���|��3�4�\In��ی��3��ŧ�H4�`��[/.u��^��̃��d��b�����m�kx=�g��M�H�����R�l�| }2��/��]�̢jʖ������̝N*M0�kgU����`-������c�=l�q,�a���Ч:+ :s�aTo%LU
(��Q4��S���8�:��&�v�2�?�<�h�'�+�U`ӨdB�;W�m��f�B�����d���A���3mIϵ��nq���e7����3�C���_�`���Ur*��� h*{���3�����H��luQ�ʬ�He�wK�S+��_W��{��m�r�o����h��=���W�(�L~>l+�Ő���ɤ'8��#���m�<�m38��c�:g�`;�0"�� G�8,l�<YX�2�� ��)â�\o�vgz�zlD���Y2���� պ�Rz��
jd�m���j��0���cf�H*&�b����7��C�J�l+1g�<�K�����L��j�����������q���!%R�u�
64][�^��PNl�?s�yX�^�w���M�-�p�wG�]��嗜w_�~ Yt��l�Px�Pr�&
���y`�e���1R��.G����I�*A�����T(h�n�þ���܉��z�l��<�\Өt��VG��k�שn"�0J��R[sk����ӘH��4^���=em��Ѥxg�6(���&��������%����� �[杞o��AP�H}#�����2�:����jLPK�7�+#:oz�~��f�4'r#�}�0���h�x�[qw��dw�5�%����L*.	��}E05���DvA��0bp��HUgn��h��׬�`��fD�Jn��z<-����Y��\-����t���A�M�؇�SG!O��֬�$7��EZ0���K2�,@w�n=-�-7�Qe��(vc��7�5��)~���|5Rn�H��\�)���2��Ex��]��h k+9����Ps���1$7�f�WX0�L�3�˖nF��xɩ�@Ll�$��n���KK�m��0y��"H�8��gx�M��(�n_!�ֹ|Wk��e��\� -��3��b	�W}7��yj���	��a�s�ыj�7�s��γ�V�HN�x�!�bR�Iyɋ�������)�"ҘrhM�O]r�X�:G�_�'�Ia�U�[��i�#{!�Yж��M��_�2K�Sa '�����l�nj4R�縺��o�"2Uz�	��l�B����)��v--��PE7.��H�w^>w֕�ړ���U�3�D��"��)U��?D���/�e0?[ռ"�=�N�YY���w����0Xٜ▃��2��
�wXL�U�w���k���+�e��]-�Ы�R/����=��I��2)h5az}�
�b�׮*s+�+m������
��ܚ.����|���,�`\�Kߏt��F�-,�1��$����{�:a@�-bv� /͠�O���{C|-�%��.�i�I@cah���V�D��I�;g�S���省/��]y��~n�T1�~�AUr
x���*8�����J�B�\.�_q�Z�k�Oz��d:��9��i�.G �w�A���s
������#:�:���Wt��������q{���'�vT�恛�б��Qo��n�,%PC)d���m�1�4�:�R��6T3�|����E�5�B�}�F^�$L0���w��ܥ�{���)��ޟg��f��:0��٩d�^Pgb�����}с?<�ņA!�ΝP��+���(AS��������5�{{�uП�y���'!R�����/��~Ĩ��a�����ʹ�p���I�ʒ�apYd(��\l�G�b����aﻹ�2
ۖ'�[/��y�����Њ�Lk��`�(��_���ϗL*��3�����4�D�̱G/��.*��Ih�h=�1@���{��Y�~�������s�2A����m�j>\髝ע>%����p�=���D�r��h���TM����v_aV9�@G��W�D�*{����G�"�	,v�Fm��ʨ�M'���oh�2+#�=�q���n�,��#B�'Q(`}+7��"��h�0q���	6iD~����Ċ]���è��#gu�oLl�H'Z�7zj�`��P�H�#w��M�֯���$+t:�l��F{�����E�=V=*�q�r0���p����3��L$����8 (��pT�����<�� Ӣ�M5������*���R?-��S+l�"T�Խ�w]E�=�aC�����<ڭ��w�U����Օ0�\�� �ٻZ��+�_e:a�'Ӟ����|����i�F�w��������Uզwq�:�(Q�,�N
�XN�"���X��K���ٙO�C����X�j@mzZl��8d�����e�q��e�����jF���+U�/��<d%�'�Me�&f�����Y=��VDU"?�cw����E|��Nw�[���{���D�2\��h:��A'�>q�GQ��?G�K�����)�����q&��8HԱn����ܭ V�Mu;�륀�*�D�?(��oQup�S��5Z��-�	���Sgs\��Z�w� .K�&�ocec��4B_�2w(���낽��l�"�ɘ����-8"|�i�4��R�e	��GT�oԓ���=�?�UI��ƩNH>����Tʴ��Ԭ8�af]����;w}�;K���2 �vT�'���̎B.0H�f�ܴ����Cd�HYqX���ñh�ꡲ~�r������"�9��]0�Y- s���°x��Wp#��,���,��K��f�2�)������\�cj6��ע��*O�̍�wt�a�!7?Q�+(n�q^�oy��
�>j
�o�P-��6����3���ީ�c�3n�ʹ��.o�LM�׵R�I�6����9�4�#f�-[W��>�Ha�Fa�/)� T� �*�!�!�[ֱ<��I�p�R��eD{u�Ц�B�F>A��|��|�t�7Ļ/@�4��xlc�U慽G�S��"D9�]S�s���KSDQY�_
����}ᗾ%Թ1ˍ�)e�s8�j��ŋ�ϵ(B5��-�k���{щdxIq���Mu��x}tX!!qr�-���)��?*r^��o�2p���X���֧����.��_0�v�5䃉C���>�V��E����䈐_^{�L�5�f%w��m���h��w}�_}1�A�
ِM� Ba^�V�l:�
�;����<�����הD����.+���,0�B�G���&���m[r,C�Fz�w�5�F^�y��9��>؊M��K�`r`�ދ߉�(�@؈����B�7�jLnY흮C@�K��O���b�*��̫5�&(�u_�)|J�QA̙�8ݹ�,5������8	�Ӭ�h���d�[f�ƀρ��åS-���u0�vB�gi+ﱳ蘸E�rcz)\mO`����XH�

��Ke"�i�D�ʁ�Z%-�'�/���,50"��9k��j���ik:�])���\X�e������g��\�+�A4@��*�,����>d���(ܚ�M���# ��C�>?����p}���nn�������wG0���-�p�B5h�-����F3�9�l���d�����P1��O��>�ˉ���	��rD��1��ʱ%�iY��aW�̜�"��}�z���U���>�����/�?��^���l����"�tJ{؂�j�����^M��>��*������:��A�J���^����΃qT�u{��=b6Q2�ն�i0xdB_���ɹ� �s�������Ad��k��V�,�y�h}W}A���' 6ȴ�=�rXF�����o�"�����MG���~ڝ���o�X��t����oW�
�rke+�^�GL.����e��*�e���N ���gk�&���V⺮٘�9�𦵧@2YY(:G�*$qQ{-���޺%*�	'�A�&��DLD���j���p>�pypEAT��ׇ�c��j�~��2�2�lף]͌�O\�k�b��X����;��������=ʼ5�� �J|uz���N+�e=���.�fȏ��s��P5[ϏJ^�\�y�a��əʖ8��G�KS��'U^^��e �V�;`fd�cZZ^�'E
��]*�q�`u���H�iD|"bd��ɤ�����8�G*�Y���	g
�JN���	�,HY-�7*�'IR#���HX�|F�\���}��l�[�ߪ"@-���`�/S)C,��/�e2�%j4de@� �k��K@l���:�l����%X�B8U'����{#���Ň^_�H��ӹ��O�v���ɰ7�3�Q{.�_$
F[�(����.��#�0�! ���v�����sk���D���aKc%wR��A0�q7W�F� ��N����@���ި����E�[Z�X��sej��n 0~e�</?����M��]�,�&�ؽ��G��rqy�w�!��h9�Z D��e�/��%b�d�57�0��hL�eG/���4���xė�u��g�x��^�fغ1�)%�ɮ^'�Q�?gi5׸z�5�˄ݓuϼ�C�:�)a��Z��}X�9���?2�p�ʈ�lc#�?��8ד�� �˯M��7I�yo"�l��g����`4EGր�Gr���A�i�隀P�ryy-C��]�����r�S��,[�z�%�|��I]�%���ϟ�+(Νg�;�j��Z�j1R��&���%�~b}h|�������;R�N�T��/�(`w�����N�c�~��i�K�:�M挰�\�L�}u�T�H�'�ڞT��Djp������.'�d�)�1tәm�A�'N��ǖ�ؼ��
���H����aV���_�ڄ����}��p�(IEJ,$s��R��1!.A����9.�OZ��+�]M��e�!A�E�}�/��*΁R�}: �K|�Q��6.��'qތ��]��P�e*�<\�=�S4ȍ��8����b�|Dٱ�x�Vߊ濽�鴤k��qb+a*cE9g|2��xmn��
Ϭkz?����Q$A����f�$���@����~!fe\���@8R3G���x��g��[�k��Sx��"�K�������QU�̓���oAj�#a/S�+�~m!�ޛQ���ha�]jt�]��\l�2�s��J��K�r}���t��_&�O�L@ZW�p��H�`0U��8��u�l)�m��""o�B��8���y�cޚ��j�J���$+�RgЁ$�;G��Ȅ�u�Ļ��2y�^[$�ST*#cT~	�u���b�W��םһqĂ�"d�R%� z4_�B� ��:�;7�e$� ��h�r�k}��9�u:8!_TᲚX���Tj�B�Eoe%�%�b�Cڹ�i��U$vT��.{�e<�𕪅;���Qh2,Tk������`K��.M
���(�����L�NBi��L�]�Y5&�@����s�)���%���B�t^+����"���cB	�	��*!l�5��t�͢*�*ٯ�i�`�<	֓Z����.��-�A�R�J���T��~4���kp{8�eV��z:Nip��*�I�G�������k��j4��J1h�)�T�Ւ�T��^��[�>w��V�a7�v��J#X�8'���J�e,,nE�9%���n�XV�����ܜ+�nFp�d�iU����A��P��"�k�a�}��
d��;ٌ�����������O)2�ǰ�OC��_� ���	�X����Q��;��e.X\����K��J�wx[�TO�������z�%�H�j���=ui�[�g��8`���u����{i�3oڭ. ��/|Mc�%�蟸� ��jP���C�AKN�6��Ɨ��ڏ2�LH԰���I/��O���{��e��)�x�T$a��72)��4n�3ę�8���_)�Rd�/x�qmZ1�-�/�n~�h�}��%+�{����E0q�hy���Ե�oL#P�B0� ńXg�L�;�J���`]���Bp���:d!�%5B��j���"����6���8��,�k�KP06�C�	��
�6@|� �k�l���G7��/�@7�{�x���z?��1\گ�Ɉ�F�p�9e�/�Ib��%a�W�9��#z)�2PD���X�R�Y�	����S���ZG�"&����\����"_�>{�K�\�׀�e�e��X�~j��h$i�����H2�%�a�1�K�E���~�%�F64F��m���ư��iR�b Ю��AD�f��w��p�.��J����2��gG>��P �Z�D���GA).S�Π��Syr�)�c(X��J��� �dt��PX����<1�>��O��<-��rߒ�"�xITa����Js�1]Wx�b��3�E��3����zK����1�X[6���4�q�����}!xSɊ,�J��J�Jo��YY-/�p=T�Ӿ�� ��R�c�U��d7䱰)<��Ҹ�0�'H�N��'~,�
�Up�u�����A�!�u#�j�g���2i<�,H9��Hu��a)1N�܆�,�7��i���#ҵ���0w�4>�t@x���/����%:y9NSV�j��G�o��!]e`0����,<�}cߍ��v�5ƨ��d:5�[���I\��ڌ�I`/�AK_^�s}�י��W�R�_b��̤2�1�A���^	�ܘ����0��|UV��̀@n�a��
/�K|�)Q�`������[KS�E�_+� �K��Mj�6����i5d�o4ct�e�ؔ�/[������;Y�#'+(x��9���֏J�4�FK�zV�|����"�
V�l���%�G���u[v-��4AA��vc�d�/������z��|#3x�
�ă!U���G��ң�9�{�'�wE5vf�;�&�K�x�a�_>F��o�ho�U�*�]�}q9�Ӯ.�<��uN
���h�_Z��]����ah����̎���e��p�6l� e7E�;�R-p�t��̜�pk}��t�a�nE����wi��oi���ii�M��XtYg�t�9�>��c_:��u�(΅N����=��(g�M.���,ͥ��^~�Eï��{y|T�eI�>A_1���:��`y�V'ZhT���[_j3F�]J�v�lB�������X
g�h�}o`W�
���`{��8(4�j�O���@���@;�zvtM>�j���r_�(Z��������E҆j�f��rg>�i�e��P�hr�����&:(�qM�e������ι�:����a5��+��#D8(���τ4Q~�0�T��e�6���ܵ��N��H��t�,������)��7��Wt���e��d�$-sȿX�bZ��4�2��ɪ_O��Cq�-!q3�Nk���&,}�@!��KҰm`���J����P�,�jc;�����rS���P:��gQ�������2�J���R�����@��� ao�u�"�����u�z�7 ��-�o�1vhG+�&��X�#�*��W.���3���c�2�}�d2�,ZN�/��u��E
%�&���
	*���K���s���� j�?���Y�\�{�Z�\2k_�*����@�m�h�Z[��Ci��=�`(�c���و�̓���x�[coWL!�E��6� �J��\!Mm>�1�s������x��2<�}1ʺ�o}��<����%�v�s��'V9����g��Q�:�v����X�F�k"@,�7�\�J���K#��!��O}Bzkkw�ި����IEkJ�>4�v��Wɗd�ܶ���ֿ��d?ɇ�ZF_w� ,�/�����n��6m�b�^5��1��^����҈g���0S�~��󝶖���[�{�z��AL�x�n�Z��rӠ)S�t�88�D�]��=y�@z=7�Ȇ���s��YFx���;�ڄ�LnP$cp5��~T#�Y @<v�AUғ�42,U����o)���E�\��oy۳�lm��~����� +���6���P��sZ���޶�B՛��*n�OM��&lk�7wdagѓ�i�ʪ\W���u�i�V=[?te{�����k?Zw&rRP�_��Ț���ǔ���ʧ:|�����b�@n�`���եk5y��wG��h�*<R��΅>����Ξ{b���;�z,4e�%G	�_w9�Ue��s��+�iȷ�GE���@��a��`I��s����M�F�-iX��������0�����7��u��Vn��Ɍw�s6��Xr�Oq[VЭ8�z�s�禰�cs�@�k	mhOJ�3�EMlL���⹒*�$�W_�7Բ��(�}�,�q��(\��	i��g�ġ͘1@`��;����C�(w��AD���A�s^�0���\!��/�@��'&���Ὺ�'�������o�F(�eU����ey�����})6�������Y�J�d��V���L<k�`Sa��A!iz1m
(�#ܼ����/���";}��[���`� �i�u>��'�^��U #_��3^����ab�2�f�䀕87���o .�@�D����N�����m��ə<]8�s#��̽������Z!�� $�q#d/�n^��wӿ���S��8'�Nb�Z��[�ؠ�O�t��Kf+��޺�&,�k(����n�_��G����'�|̌�P8���A#��Կ�#?9wnQ�ܥ�H���5����0�I$��߫݁ځ��d�eW7�t���^G�)��^�F�����=�Uꋲ5mX�fqP)�K]���7az�㱠/��B��v'4g����x
n;�ǫ�T�5d��Lw4������;E�[rB��bJ� ��m�6��67E5 �<R��ßx�|�e�����t@#S��5}���SՇ�y=E�GzEv�|��N	�L�?����H�/r#���-��r��ɵg7���
�_ߛ���[⓶_v�{�ٵ�����%w5{2ܛ`�o����H��&� �e�a�[6�p�w�'ƪI�@d+pg��+���K*�߇�/4����c����3x���������ȴ5��D�.�=s�Yd�*�h"�#�FJ��v��p�P�F&B��p����8θV�2�D$Ve«����z/�F|��dH�C�
V�
��:B�!cp���-�N����)��E�`�Do�A���M�Yj��j��CCW]���!�F�g�m���f>13J���h��;9�'uO2X-��[6S�A����LZ�K���ű:��5��-�����Q�[��#���DC�^I+M�C�esWCr��Dđ�N�Η���<
iҌJ�t��x?"��t��m �'�j\�R��E�B��B<)n��ӑ�
*�A�\�h� �޿f����`rw.=���H���=P"�t��L�U>���J�|�C7��_�zǖ�n�+�Nhf����Ȃ� 9�y>�sޮ�K�����)�u� =rhÉ�	�G� ���_�B3�I� |�T��8D}��h�O.�Ԉ�N�n���@�->��lLG�<7fR�Y��� e�}@G�V�z�3�(.��'
�T��0ہ�R���x�k��6����)E	;���lv`���^���HWd�����q�Ɏ�5�٪���	�I+!4��τ貮B#ӎ3*ΚVR�]���=���I݋�7�\��?���$c��-�@�������m��7��-��(ۙYgM^�%��2f)��3}N3rB�.ۢ(�J�.��*��������1a:����4����[����>�RS<nT���N��a`d�$�pxH}�Qs[����Y?�20����ְ{�EX�0';FN<�D����&�`c�lX�]`�����e$������g����8F���{������w�)� ��R�Q�y-2�	
}3q���t�!X���a�L���ۅ�Өؑ���gvR����ٱ��k&_��~��$u���\�w�ߌ����8@|̉�:5?��ٗp�D�߰]����iq�%�^)�8Op����;oA�|�$��!ʣΐ`Q�|�u��e��b�I[U��%��;��\�{��]{�����qVF;�:��������;󽀁�Ӫ|1}�Jł�5�������H�*��9Pj�t�|%|����N@�B�0���"S���\�}���M6�)���Cq$��@�� �;��I/jtq�c2)y�Þ8�|U8b#�+��T�z�=�Q�h��8-h��:j.��	7ک�.nχ���1B�a�x�w���5��ΜwrQ�	�lD��*�ƹ丂b�bX���~���2�~w�K-�\M�	;y2��.F�:v����� ��i�MI�?E�	nv�QiQ4;u噭m�*�/��ѱ�:�\����]�>����4/e[ǖ�c�`��d��	�����n�$�HK0B@ ��4�5"��,�oRUs�>i�0��kD0��Y0 �HSw2����O�+�n�y�wH��
�`�m���:1����ɠܳc�l;��W�?�)��L)��^LM�p��Ey��'Q��q4�Z�g�ʳw#f��e{�@�L�����m還�J��г�@�R�e��'�kJc�羚�ݰB����=��`�9,ڑ��$�8�Z���ےp��s!�M���y�z��M9ꢃQ55��v�F������V���¹[Ƌm7a��^�~��ak\!�DP~�}n��M]��o�C����9�L�+~,J�*Ȑi�ݦa��6��]f���M�������$>�ɾ��{���>p�y��i��ʜ�.ML�R%_<�����֭1�܁���S
�8D��iU�$�\ô�q��P�}S�B^K"������01c j3==��\n���e2���Id��E�e���Cn���/������dw��#)��"N��-��0�����y�� ���]@Y܈�-��!E ��G+Y�#7f��S��I�7�ϵ|S-&$;j�u`��q�4]����v<���9
'���N$c�� �p�`��)qQ��GFm��UW�h ��e�4�����CۇN���O�o��F���G$\x�*g�~�*��a�41b�Τ�kv/[��ϭ�2�����������+��"�=t��D^&X�i��I}1�a2ҏ�H,��K�4�z����vZU�Ud���w򆖺lSn\��s
=�w1�@?d�Y@u�O���5�6z7��Nj�grˈ�CI���ݚ�0��� X �-4��[���fu��@����d��P[�7Ts�G~"Ka�?����=>A(���4�%��A,���]��?9�"e�8^h���6;��&�V^t�S�g�:� h5�ĭ� �8Jh�C�G���^��?(h?.�ˠ0�e�=L�h��|��J�',���3?��gb���841��u��{)�)���ԫ��Wr'������62%���!�vF4U�������;���Q{��GX�)��RZv@juW������9[gi�"J��8�j�9oΫ��5�cpq<ttO:̣&��q�H�K5y�e�ɡ[K��.mn��#�_������ ���ɫKV"5KN[��� CQU�?���I���12Lc��C�D��h���9�c[����6��"��Hr���t��j-��-������kZ83��Bj�7�湢I���_�]�o��/.�U~c$���Ch�����K
8���a`�3�O�wG蠁T�����j�R���"�9̓��ß��$m��	Jr!{�+8���F�Z�agzX��B����{��h� �6P��7Q�x����%R�?�Q���~z�[�|�E��_Ai�C�1�1���<���.�� �6*b/K�ף� �a�0U6"��� ��8]��"����ED���/wA��*�����Y���`�6"�hΘ�:UwS�s����A�C�QB,��%dNH˙�ط�F�j3n`�]�4~�`�!��k�k��˱�'�;(�V���q2�١�T��'l	Fuv����FF�f2U����Ku-�C0�"������1!a|�n\�RK!�};\�=m~�~çd�����SK��ܚp��5�3�����c�dkQ�zT��-�O��`��"s�K�� lS��J���Sy G:�
��n����J��Z�Mmw�z�dt��^���Ԯ�����M��E�@�hT<��	���V���'����,���X)�@_к�IE$u���}Y�MFQ�`V���3C��_�	6i[B�d�� �b��/.����������Y���8��0=qK�k�'[�I�O'!S��m�'oD	�%������L�W⥍����s�?��9$�6���Տ�}��0��	e���8�9C�pl�md��a=M{n@�)Hq��aǔH�������)Y�9�<v�h���G��c�M2[J��3���ʃ�7�@�LBs�dr4�΄�eb+��0��!��3MǦy�?f�ve@�r�/%� ��c:� @t��F�0�X�� �L� �ⳛ���n�V^����nM&���h�y�f���l�_���J�}�̝Xv@�B]�P�=_��ݒ˞1�\�����]��Q����)�)t4��Xn�:�>���-�x�&��]s�U=j�һ�|�NƓe�H����?f��jc=�ը�^�  �D�t�wS����I0���:W�t���,��ۆ�O,t�'&����%R��AQ�&d� 3�����@I<z�(��A��C�` �f�j�դ�ݟ�J���~�@��23L���c��W�5��_Gxy��WO�ؠد�%�[G��?<�L�R������&�Ƅ ����ؘG&��{��뷰���"w�+
r�բ�x�\��:��Cl�m���ON:�[��
��������70�!��h��a�96=��~��e����2K��Ì,�Đ}~_��FcSZ����5�$g����;�/〪����HGQO��w�|��s�Y���\@市oMoQ��ؒsA�w��r��(��I��~(/�_>�3+i�D$�6���u�9��`e���OO{┭�Jw�:������W��I�=I+���>4f^vu=�[!�Q����q����T����8�� һ�٨2 ��E������Q����n:�ܲ���`�8a{�&�1��J-�_[�p\�ଠh�e�!P:�0��+���;���v�
w��"��wq
/s��E�țߵ�4E��d?��c*�,"ijT"���:��=��KUb�K�"AR�-�y�sX�T����֖,b��'���J@�Tܜx�A��Z���W}�(�r�)��v��z���);޷�;��I,6�:,M]R�ں�b�X,�X#JRK�(r�K���{��𫼌��6C��ͱNK�������/��~~���b1Q�}����E��GE0a�wJ,�:�����sN֩b�hұe}� �y�lY]	���x!�w9k�lNषW3�ߧ�UX�F������_2LήTKڼ�;�M�Z� !��нoc,R�w���
4�
k��������K�'�����V�dJ��Vn~�	�~�;s��ǥ��O� �B�e+�%�E�����95z�A<��т�o���ob� 3��st)eC4;�Q��z���b�RVrn�ڳ�Y8�+���6/:8J���w|��\�-�Ib��U�Tm7�[�$g����p��tо�Ix��8N�)� �ٿ�94��n02*ÔK��)�"���݁E6��k�y���y$<�L��yX�����=���7�c�LP�X�L�)�������Âd�C<��*#�%Ô&a	��\y�,����a�s�59qy�b�>���Mw�����b-j�?jYXE��i,�o�[q������ն���E!q�sj�v�b0�?�PeY,	W&�E#�u���H�W}��gFС0o�l#L�.��!޹��2�'���;
�š�9j���%7=̻ͦ�[z�UC.2�g��o�Am����ĭ�5��?�L���0���?!��ji����o[q���%�Nҝ�Q�8�y!�7Y�����C�[6SW x�W��V�=�~������e���V��:�Bc[��{5�:���z�_/�Y�8�\E}�Y��54E���t)ui�+u|/��>�*�%� �9�`)���cc��#�[��o����� 8Â%�)X��Sw��)�Qi��k�l^j�X�x �:v�� �!�_	JiE8~�|	�3�\�4���ޣ�ڲ��[Ob�4�k|��ԁ�i@rڿ��c2�,����"Q5�����/)� E5���:@�q��LBjpE�r�1���o5��X����`��8���8�[���=Z]�s�1>lO��Q���
��A�ŕ��ۀ�>f�g�����9� �Ĵ�$g,ґ:���0�(���^�����i�})MK"gfHZ�xYY[ͷ��9�u4��6��.���]��耟��z�:��`[����S���2"��h��-i������c"T��/��O�K)n��Zi�L�~���}�����W�^�
�7ߑ�ӷ��x4U�ս���( �ﾑ�����ao��� �XŢ(2p2�`;(��F���2-��޽L��������S.=1������D2�Gt��)μ)>A,���S_����{���A�E��޶�T�2�P���f#4�E�9K9Y�J.u�e/����$�	6�%�_�������ys�r�������F^��Y����х�#������������H[�]V�����{O=3��@O{�i�2�V1�xw�a�{�JpHu�4�u8S����,9�		2\�m&S�y!����
i|������V� mm��k������\P�G�Җ����+"�(W�mj�du��l�;���?�t8q���g.	2��A9��M�a�I�d���F�ҁ�v��N�΀V-�$�>���2f�8tW�}*u�\�%�{} �ǌ,�����)���}�����6�YG�����S����j�v=v��OY�H�0��8��,����
vpN��(�!,)��8mM�
*8*,�k��D��������۞*�&��;�/%�m�[�ґH���tR�$9Qb����}�&妯��]�Y�)�#��i�?x_��B��<���\���� �K�0��*f`xo%TLK!�˶ɜ�	W���ՅqF0�N4X�w����Xa��R\����z��Ⓔh�nh Tlp��չڛ�e���v��yiK���8�B�*oV8-*����L5>��	�2����'�U"�a��
n��e�E��%f���1��c�[��NT]4 �˹��ƬJ߿�+��j��vq�~80z�5)�T�X��0�
��sU%�٪� ��7����.�6K�^	2����FW �Ύ�����heAr�י�&���5�]�	͚�1s1;���8e*��J�bƚK�N86�6��}D�&V&YM{��b��\�b%