��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����>�S��fI#�l7x%���$or�#�6�y���N�i� �D��f(�:eǊ�` ��S���^�mBƱYjA���v�0��kh������#�v�(#W��ux��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htdʮz_�0�`��@�[D˂8��k�ľF�n�Ԥ��r�τ�u�&&����\l&�$������<H�����}�ƌRS>�(B-~�� ��ڣ�9#M��c��&��C:��pǾE(
'�|�7���UE8�Æ𚮙��U�
�'�����5�:c�E>���t�D�n���j8�u.(�hX5'�������4��O���vݦ�Z�Ğ �,�#|��X��~���ҭuH9H(kk���)l���m<Z�� �ٙ�N^θ*)w"�Ju�7��@����a�nK.���|�Bs	�o��s�Z��q��z�4�D ��er���iai�z��D��WO��\xO���c�����:�����T�)�w�l�����p��t���O�A��@���_Ky�YB�y��p*Zz�|c��	�ٔ���DT����O�r������q
�&�pX��"9�Y��4��E��f�_V���yBa�Oo���vu��Uo�����c��8�/m�2��2�y�ԍ�Y�,�Ɂ�/:.}�ӊ���*�C�C�J�<e |$U6�z[gV�.;;�I�e��L"	�.'ү�!0��*���R����3Wf��J�2���ת���smrr�(5�TQ�����Y��rK�>�u$u,��/�����W���q��w3έQ��n�\~d'��}4G.!�㏂`���=wq�@��I�ta_A:V�>D�C�sQ��Ϸa�7U{�P�������=�x8�%�ff�ʽ�Y�q��e p��8<~�/�����~%vSuYOW$�MJ�U����|z�u$e�F/����ۃ�����D��SS�o;¤�.S��_=�4�d|��X%��n�Ɏ��?ӭP����t�x?�|�.F����C՘��t����I����Ȳ���g5�wI���p��`Yx���x~���5,s��Cz`�l��w�|�E'C	2SKt�����:b���~b��İ�E�7~�OZK~�島���K�vHb}q�t;lԥ��-ʰ���n���e	��Wm$$�ټyͺ2_{�)�ȷ��#(6�*ԉw�)�gU��b�<��V�%�;���u��i�P�< �KZ���VI�[5��t%�X�%B�(5r��;§(�؇�I��Zѓ��f�!\^�YD���_YF���i���D����'Jl+��`�;k�	O�}՝QN	?:E��@l[�Z�s��i{�X�B��90ؐ���ҺBz"H�ef�<{�pr��8an�ݳ��H%�?_����u5�?��>��5�\%[W�j��T�c�	a��
h�8
Lô�Z(���./�c�\)����U��_��I�t�^0)Z�W��v	���Q]/��s&�/�C������j�$����Y��W7�c}�)\̛���$��#|�nK�����7WE��ъ��������D�6�^��QνnFFS�b�c�j����sy�=�I�I���mb����O=��=��y��<x"���cp{I9��t���^00�ؿ:�s�FZ)�\R���k� ��S��}�8u���q�<peŏ�n�;�^���_�J���#?��������r��:v�[nW/	��&|Ml�kÑ:p[O�2���NP�2�*��咪݌�4tS'X�*�|�A��Fe� K���)��7��Z_'�N��� ��d>66��{�-
���h؏�`,�AS���t���z��Dw:���8p�-���do���$Ё=t�?i����&ƏS	������0mZ�ষ�+�Cn� OW/��K5�R�b��6������;�o�m����J,�c�Qq�SعB9ʬ6	���-���.�z����X�Ou]�\a����u���@��CD�^Wd{�s�G��#���%ln��!�y��d���z;- ��ю@b�m)�v��sD,�Hg@�hs"�
�Wg��wQ5����gUI��(x���!TF)�>��=3���|�K��;מ�Ň_}�1W�F]"����;���[D�D���@)�U�'�$n�������X�x
��y������H&~z�GB�I�2݄�g�d���r���B1�L�c9��E��/K����Z�"��(Pkv �Ż�"�a�$m&�������z��2����$H'�5�n%����p```b��}3�%)�"�з�_ ��I�}�J�7�%`\J�KƁWX��E�d���#��No�h������Rg,�����Y����ٴ��T ,�6�~w��|����n:I6h���?�Lƶj[�C�vDT�����ǑX�W��,��Gs*K��,>�
F^°��1P�D��e�.!(-o���<z��������n:oS�.��Y�HQ[K��2S�L�-���w'�䞈�k:���;H�!������D�@r%�AV�NsJB��m����W���m���r��|dQ��5	6O_��|������i@ut����<����,?�G�ߪ��JY�#���Kz�_��?��#D)��&�? %�w�(v�P�'��N2��V��^���à�<��,���iZ��|�c3�Ag2��x�����ݠM��hV%�*���32q)�W4@g�9;F��|B�N�<!=|��_v��]���d��hʹ�% ͉P0a$A���0S��H���������C{Kuzr)�]��������u`��6���U+z���~o ��+f,Ǝ9h�\c��
^�woU����(}���P�w��%ZC�!�P��1�o�����y�t6a����� �k��������օ�5uShu+S-
�x�0)Y��a?��疿WP^��̯Jg�V��&���'i�r��J�T����_�8��\S�O'bֲ�+������I��K���#*L��
��w��͜�ػ�	ge]��[�7RA�,��et�_4���:~��gVU;!���7�'��ǂ� 9��sro�ML �h�V�ΰ9��xo�m-1S�'�{^LF��dT.�2�6�p�%C[y�$�J`�K��8C��vѧ��F?f	����E����ccU`����Ls�6���,X�ۦ�:���Q���jL�l��sml>X{�����]g�L��&2�d�.�'�}>-��vs����a� �j�l����`�6)�� j�x=���,��>�޹tɀ�d/�Kl��e�\l���#��ņ"�H҆��o�I	g�g��bU��}��a�g�VU�&�!'��;����g�Z��R��M=�X