��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����>�S��fI#�l7x%���$or�#�6�y���N�i� �D��f(�:eǊ�` ��S���^�mBƱYjA���v�0��kh������#�v�(#W��ux��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv ��i��X��s�-�Q?F�`Y�������� I֏�׋������H[��9����ۍ: ؕ��6ж���Q��" ��y&���Y	6_���.���M�ݟ����k����
۷j	���`a�s�Yot1H���\tr	��:o�88��5���w^H_�.���~y�o�ض�d����_W����K�3+4��-����0pl2<�8�_��%�W�!����5�#�kͽ0�Ťq5I�Pkc��|��k��h�6���3/��c!�)rJ_�t�$o��1�V��tGH��#?��a b�gYG�>[��;&��Z�M7w��x�΂��^���x�*u2X	���+^@�.���;�v��^`@)^J;�Y��O��/�������8��[Zۏ�[�%N/�BAJ�՗;����י�$�q�h���%7ev�x�;��GM�ٯd-�������!�	%�vę橷� �ݐ�ZNR��l�Ȓ�����(3�@������#j�7����-Q_�˺�wZJM������*h�f}`�'"�3fM�k��ys��d�?j<�wB�,��BU;LT%�k/0~=�
nP!��s�:�c��l>&B���֑�5����se��W�I:��R�1a��N[Ng�&�W�7��ry�a��S�o��И���:�-��?�f{����-�ݕuW��VD��Ke@��9t~X]�q��Ɇ�uSQ��V�^�<`�n���Ҩ�h��J�S|�*fA�<~K`��<�Q�l/ ��KIX�����=O��w�	`Z�[��B�U.OY��PT2F{�H �l��Z��L��H�NߞK�ߔ<��^��gk��k���o��`�ʃ�Ir��)էUt�,}&0�Ǻ��pF���Xk�OlTJv�Lr�C�� '�m�����th �W'2;�~ý������FuQْ����$�=���/�����MS���<+4It͂n���rܘBX/����~�<��O�9Gh�X�%�_D��5 ���')^�E�!�d%	�u4�mb��(�����[��1���[7W@�%؊o��p��^���)#js1��fJ[��)�N��Ѐ���)KY�<��Ri6djkl*-���1�%�ƥ����OQNv��fuIZM�#�8w��!� �c��bP�ޒJts�Z�+/!���	j$7�6	ZrCp7�ƒ3w�Q���b�����Ճ����ߛ��x���1=#�* XT���*�t�����,㷩[�t��{y��ً����+b;T��A������C�t�֑b��7W�%$�bI����g6�(B"����Q%�Pm�;��m��T�����e"gk/��Jxa�cQm�g�WI����+�4���=�YVl��AҪ+o!��'&d�|���TԺh�Y�x����[�*:뢲�}q���(��c(v�g8憕z����;�z�MPZ;���DG�?�jMW_<J��D�a�162=�g�[#g������^�P�[�߀ݸ�6�����\���]��H��(,�^5�?u���{,=[��ṀOf�?#׳g9��us7G?̵��y��o_�3+%i������I^�?���tlf0��}L�(��y�'����
��9^t��d������}��ST�GNL�"6z���� ����|k���Vn;�E[�� ����CL(]�9�@!��Zְ"�ɡ:������+�j��Nڒ�G\jt&3q�z��|J5u�t��$��^"��h6�}m&vaL�6w�|��_�rGg��'rG�G�Q`\�Y�Cb��.7/�Ո��̀��6����N!{�KW���?��Y�zG�ǋA:��Zq����f��y$��#���ЋI����l������Xn���V��K��/����hl9J�]�x��5[��W��?�X'M�2�2��%%����r>��WX���~]�����~��-�,�J0��V��H�x��à�$]F~ԑ�����1I�0��OnG��C[?�y����|��op-"5`@��ӏ���;NQw�Vxe�b�݇s|�L��r��!8����A3�*��n�2������A�o�_�̊���΁�NRɅD<��x�g�%�����Hv�-\�o��6���0WBϹ$Q��k���T_��^�$4��X޻��_hvs�
=鯄�Wv�"�GU)#P�Bݩ�b�b�y����@���f3ӭ�W����x��
�`�8�hgu�;ӀC�&��l�]�sAk���t���g�Zd�f��B1����/����*��b�ʡ��nϠ�);�cܮ�8��{��W����Bl�#�3�j�.*��f@Y�j��r�Gf�HuG_�s����Q��p\SYiOp@�A4� �]����ش��z8���$x ����
����U�[/��
 /��ᭃN�G/��G:K��{�r��GQ(�̓�}���V�{��.j�q��ĺ��f=����\���tA����&(��rq,���(������Nͨ�����p�M(I���1`��Rq�����"��,ⱸ���t��]���Ӊ/���Zwh��"Z��c�iJuE5k�AP�&��>g�C�;�Y�ϙ����@��ߺ�ii�MV^Sm$�^��O%J$��0%	��/ J�l$CP�pP|P�ݖ��{8kD�	���Ω�λ���6�!��J�����~�1�[���ђ���D�9os��߁��pI�SF�Fn4��ԍ}�k��#͞�nJA��W��u���o� ��N.��Z�f�<����ⷑ�=��p]є��2�	"צl�ī�֯@VbQ�*��#Up��nV�=�l����0Ώ�0w�]~Q!rښ��(��m�&�����@e�׭��L{����s�O�����oG�� �AdM�������=k}���a�H�65��p��zv��eSUH�T�^�;�c�5��*�Yaf��XCH�1	�3���QB��@�?,^�P$�g��jN �t$�%���Ѥ��6$E� �3�C)��:sP������l��Uo8-�+s����Js�� xV6�d����FEW�%nֶ��,+�BR#�n&v+�b� %�}G����[�nj<l,,3�����)��'=���ZU�F8q��5�)�^N�l��ׯ���N2�����`K��f1�P�tM������S�"�Q�s��P��y��E]Á�uf�C�N-9Q�g�Qs��ҵ�po�Tf���Ty��h�z�zu;����Yk��W�o�0��,+��2�i� �B�F1�t������U��N�'	a@�o��i�ʃ4���p��[��%L0�]�8��Э6��a�<�gG(��H�8I��Ixe�Y��A;�����7�~r~
^5?���X7/�o�6�ʧGV*|џ�^U�e�K�xt?>�-�Q�i1�i�y�u|��� ip�+�MTw4����c~�%�%G$R��z�CL-�	�r�Υk�0
�R��EG��ٰ3�wI�e���F�e�*Б���j�rU[?�Y56��2��A�8S⚧�^����d�swg���T{�t��l�3���|_
���S�$d�nG�s���K��^�ի��BE�5���*co�J�u���m�����ߒ�R�W��C�@\�E��fN�Bϝ6�Ջ��
+RxB���)ܛ?S<.o��O�)�<�+�1��\p[�g��8fC��j��p�����I:���߉�U��t%�Z��i��8��a!��묃��ͧ���'�:�E�2Fw�p�b�!��4��Υ�j������c9-$�=͇1��%#�@>5�V�ʋΜv��q�p�C|m�<�$�aą���+X�%�D���.�I~4��/���X�%.Y.�p��d1�fr���vhww�GOp7�+���x>jh*9���~�5Q�س��Ñ���D�58�djm�V�c����͏���E�eXd�8Q+��������Ij�p��U0Z�2��e�t�p��Hh��Ā-�I�ys�6� �Bϋ�3���me�����7���u�T:�j+m����j�Ή1�������y�Kޠ�pC���j�7M�ѿ��R�š�k��H�g�^�m߂V�$����	����x?����p�������g�3����`�J;a�e�w�<S�.suy�]׊t��xi[({�ƻ��8y��^���8��"�����:� �n�$t���q��})[F����� -�S:$����Ն�j����7b�q����_pZ3k�D�C��Зۑ��Qc��S���0/�E=�L/���{�Bs�F\,�F��f�1ۡ�߈q9��e�mm�Eq�G��(���Y&=%��q�(a\��/>�-��3V_��Z�wcI�5g �P�͟F;�>+*���i�`�@�8���as�rG~Kϳ�fx�Q�d����n�%l���t2�o��f�x�h�h�H�x\���#��p�m�h�恎�C?'	��m��_�.0X���9{?:�p6d$��v;ehv|i�)">x�3qH���@����O�ur�u�������~S�#I��qv&������{�]*ߦj�\�n%�.�Tj�����-`�~�%6��i�2##�c��g���LvC�ܣI���f	v��Ҫ<e,�s�,��� F����8�.(�Ov����{0��k�3�*<��xj������|�}���㩢^cQ�|�o:|����lz�����W��5�ț�_:�vu1lU����+*GC���٧��tz�t���$[�	e���bgk~�YES�T��� ���̓2e��a���X-3���
>(:$����zϸ�M�������;lѷ�L+��Y�a����n�E��Yv���;C0�$#��Τ�-��Է��:'y�&���ݧ{{��'��h6U8!:�~��>TD�*�ɤo��Ŵ�.�'V$]AB�}�����'a	6��z�X�sz��L8�'���#g�˦g�u��w��C���geͩ��«��;�_�]�%�l����`�6�������2��� �;�8H>a��<��.y0K��y��*��a�߂��돤ZAa�-`cf����n�^]�!��H?�N$��t�%ené���B���yv��n\�"�f������v ჽY�Ͳ�[��%,����V]8a4'/EHʇ`^)�]a���0��A��8W�b�J4VE+��Nd�~�P�j7a�5���hwt2��Rw���
�¥��ݳd��m<�e8m�D�Q8�'l�|Y��u�#�����{�� t.ɰ�Ok��$&4fG�Ő����Sva�}@���;Nָ��nCstљe-9�����;�@�E3����;�;�C^O����ެ��~q���un���n���#��g��T�ճ3,�{��7�w�!k�!S[��v�װ
����zwR����V��G�/mdJ��Y*���y�u���-�Y"Pút��ʎ�Gc
^�v��B�&�ȍ�ͬ�eMF���ܼjޮqc,&�Ju�C��Z�yڰ(�ʌ�9a�Sj���@b�_J{т�?N��m.kf�xA��\	���(W�
�-���wi:%�m�"P�y����bi�˔A�� 9^�˶~}Aǋp?���mCT�t�j8����ZҲ���G����+7�=�t��?�������073���З�r����؞P��6{�&E���tz��)�������=x�����*�K��]����eg��"Aq�u�!�1$����y���ސ9H/n�ɒ,�$>�ֲS�����a<Lצm��.�����2���Z��=J-;T����7m:�n �B�)0��J
Y$��V�!�*b�A�T��L*Q��4ݑ�qTĻ�qˍʒ�����\�!+�q:&��x!-/k~�*�	iД���7޾�ʒh 0UD`K����-5��#�M�sx�9/:���k2��ր�>�m�Y�����m=�e�>�g�v��6�4�;�߈�:�`b����27aV�K�b����[���1ʆ\b�>�!"�N�M���i]b�{6�b`k��?<q����_�m܄d����o��5]�M�\�;G����-���
D&��Ĥ�Z�tR�ݤ�1�)#��Hsb�zJT�Mw�#?u=��6�맞�O?�胫?
T�8�(t�]SrҴ�K�k���ř��v9?,�g�D���t*o��+hS7���s��{�J��t@�n`R�X���$����~!S[s��!Ԟ���ڹ�k���9`�@������H�H��pI,��
��:Zg��8x�3ɕ�n;7.b�~�W�x��A�F�����>���kC�1�����7-%��=I�c]r�r��{�lt��k���y
u�TH��և��:��X���/�hQE=�6��vXE�����S��7�%�a+�jx\�w���'���Ζ#�>V�4��_h�e��8p�`I�L.�kx{k��7�W�㗃�E-��/��H	e�����FJ�UbHv#��ٕR%Pp1� Ⲻ��?3��n��2M�� �)Ag��ۖh=?B4K�d)��>-��4�M���i|!Yw����L{/@<�7س\EݮX»�K�-�k[����%r+�d��L��6Q�����9�l��m��ӯ������OZ�
�!Z��v(65�L�*����3�ԐAf���PKv�Q�����N�m'�}�G��[<��4��]6Rt��D_a�b�~u��j�ba|Rܫ�.�4iBK����?�B���6��B�Ƹ�Ҍo��h�g�Q�'�P��v�+37^p�~�ȃ�7�K��:���HD�]��i ���t)�R�s�8�^�T��<�|�{dwX0;#l���E�|9�G��g��&7=[K|'r����-͆
ҏ��~$�i�=�6��� �����-����#��5}`����m�Ʋ�di���q�s��z��y�I�}�E R�=���,us�}�2o����y�?h/a{�g��kU]�q$$$:�Ɯ9˚{��ShǆµJ�5]��Fhv�\?=�v7suhXׁ�K��l�Z��%�Ù=���-|7ۑ�^�L����l.�9b�ϥ���Cާ��ʌ���
�'BMJ����s1�����-�,'J˱mS��'(4��i9�/s6����0�r,��F$�}.{�!F�H9i3�2���@�m���R�>�>F3�9J���c�YĪ�0��+���j����"^�>�|si�).�	��~�����C9c�F����KP�.��ď*��Ѧ?N;^�;���4^��8c��Ce�;n�w]nH�'��T��31w�F(�#f#c�O��ג�%!I]�'�VV�?��DT�UFcռ/���kF�n��O�l��)7S��MM�N�t>,6���5p�o�mt��=}ɘ}��V-`�`����z�>�;��^O�+��H*]�v���a}���$�4k���.��'��jމ嫺U]��
T�Yr0���	�>9�ow�L���m����(a9�,�"떎7���*���}g�X��X+;�?h*s㛹��h�,L���E|t�����3��3����W�e�Γ�(��;�)�/�5j�<%�mL 4�G����scGkp�u�ry�^Ǐ�h��q=��I��ԡ �9�D�rm9��K~=A9B��v���gՕ=�ا_����:-�����[W6&r�-ݍ�L!!;-T|ה1��C3����ؗ�Z}At��3i��\���e�/�]cYRZۄ�;~k�J� �{�S?U�4$wf�۔�}"53�����[�o�sw�2c���!핤V�I�
��E�Y� n���U8�Y�GqR��������&1
�̈t0ѻ��s�j�h��Ⱦ�߂�%/ܲ�E�S�~q���7Sy  O�6�������1E�������;���+��m��N���Gq��aJo�[�ئ�]����Ib��=r�sh�"d�t�>�g�f�p^�
�BnT ����=|7ޓ�d�S.�EL�x&������H�3ԅ���ٞ�F�x��;� @�ق|z=���P�ԞL�P�iO#6_`&�����޳�j0������\�zڡʥ��4[w��"yuq�iS�_�ֲ@G�V�z�+N����e�Z}*&�2A����fd&�;�)��ȳn��r{���y�FNXܛ{q��d�RiX�HYOO�^�c��d-��R��5��`�l�<��6�z��_?7�n��n��G��� ��a:$=rEJ._%s�[���3m���kI�u�xv����4?��Z~�+���"x�K��/��o�"&
�t�h(
9�ef͌̿@\ڈd�ۘ���~�bUǣ1x5`}J��Q*S�C��7@����GbÑ�ѥRZ�_������F��\-�����_��d;Q2-ƿ>�򛌏w�M&�e�]-�����N�0 �tA�gC�)�\٫Q��ȼO:%E��A�RH�Q=�y��E+P�w�y k~�����r�N�[d�� De�Veǚd���ػ2ۂ���Й"�@��K��m�*��֕;�����&��*'U����ʂh���/�RnGN{��VuA�
P�T�l�M��O4y��Է;˜�z#kU�)�4q��L��W��1�ґ�y��Թ�o;��ƭ��r�eo;����=<�r1-Nb/�
���>橧�;�ȧ[C�����i>�����DP��( Th�>>ND���E�4�4z��N��P����C3�˄;����Q��<ҳ $�o��=��s��HK+��4\�t�r����bh��j�>k�r�q&	Wol�"���M�\��>ޓLK��M�0��Gy�@A�2�����>�p�X0�'�m/ۖse�v���ݳ��ã�޽=�l8x�||��1]�j��~n�L2$�^���Qbea�BK�	��LOI*���K;�\S�hV^pA�<U���k<�l7����!9������R�J]d��?
�`0q5�7
<��uRUK�"�N�Ǩ�t��X���	�]�X�Lnx1�n�2����A}r?G�~K�4뒵�x�Ӿ�F�� �X*� &4������I��?#O439֓!�0Y6n$�P6TabFG�&���C4�$sޮT�+#Gkߊ+����䞃e��@�s��FD��E�_[&���҈�{��[vK'U���I4�9�8Ԧ��maσ�Zl ��2�"<s#��|�Y��c=	���eV���Q�(����ˍ�?����$�M������稨���ħ�{phK�a�-5%~�%�&�����cIhݪϨEl2���LزWa�z2^7L�9����c��4�n-�Ƕ�r� ��B!;��I��Ϻ�L���v�xWv�htmބO���s��� �Ӝ��mX?+���h��q׏\=�3�{*p;��ҭ:˽k�f%��P�����_ؐH�-��mYB?��	/ƁچGZR�a���1��R��`���v���tn�L�#-DB���X�����%T�q�Za���s�e}������ul�$8pZ���d���Tߟ7��ݥ� ���U�4�V''UI�clY����xs�IĊ{��X��#����@
�-����<������۵�k��V0y?�D��j'�:��9�_�T�;}�~�n�h���}#�u�b�T��O *�#E�K��(��v9�Fc��vhB�L��o�ͻݙx��!S��T2�$V�H�3�.5�#�w?yp�F*����m}1�.�IJ��4E�[7(��?���_�f��v�}M�f��+"��5�j�S(�8�9/p�pD�}a�Ϳ
�n���|�����l��p�$����/X��U�I��Jo�,���	��5��[��*-1q�ە���%?�z57�{�o��Z_1�3>�O��ݔ���	'�2�� ��h(��)�7�͸lheU>�	�" �z�w];WX_��	� ��"��5JD��U�@��<��l�m�a�~R�gJ��h� ����*.��f�F�R��4	�b��}4�֦%��s;�ĥ�H|��j��֪i�����V�cp�⵹w���%/i��+3����ȶ\K2�l(�v���ӳwx
�[�#�ǉ���,�}��:��h�dKsy\7ƑӍ!�[1N�~L$���im��Y,��׵��9Gx���M�}^e�i�մ�vu�a��?ᅶ��FKO�Wu_']`M����7�-C�<�(x6��3�2}g�G,���c�d VmF�v�'��DT12[_"&�l�sI�,'�a�0� �R$m��uv%��~�{H �1��?�2�}�#�g}A���+��~�Q�AJ��B=E���)/�:�_�����%A�f�-��=���?�H}�6��Y};�ƀ�;��b0n����p���! {�����76�C��[�!`�j�����}8s�����X�x���T�:��,RN����B[+O��%��� p�� ��<3�K�s�R��e�������j٠�禆o/4�p�D�88F��,h�,h;�p��}('M�>A��V��׼�j�_��B�XↀWN7w8�'n�Dv�[�ntߙ�=��Ҫ89mG��yS��&��,�\�'�^�Q�wd���ҽ��t �{�`�?Q�v�l���i�x2���E��D�H�!Z~�s�,uЀ���h<v���F=KJ���p>���fOQ?�e�#�f�=��mI0�s3U�R�P�s� L��p;l:O���ƭf�� "U�}�����\�!v��&����ֱ�����;ˣ:��T��Q�M�$�Є0�V���<���n%�ف�����6�y��.��([	�+��f3u�!1ul�~�4�Dm?ty�?x(7�,TT� �2%Nf��W�8Vf�HƲ�"�_�s�2��-��˞S�1��D)��>��l�����Q#��.{�3]Ó�B;��B��gt�p�<|(cw�����ND��k�Pg�����?�\vS�<�t�T������b���G�y#q���W�W0B\��� ]�5_a�u�(�je�H:U #�~�e`,p-�\G�����Vk��$Ė[{���p+++�Roco�9��7��vɠ�᱈�+٨*���Gw��~u����SH`�{�,��9������ѷ��&TMO|eKjF�F�	��!)�2�_CD���h�{�I Z6Q:"�l��o�d��������|�&�e��|�"h�0Q��m�����:j��7wt��$�:sb�;S�eL�c��Ϡ��ϘW�����x����8��%�"$9ZU�y?�!��+��D�MI�q��,)���*{�|Å��������#/�sE+�Pv��|���4���A�۷ǈ��\�u؆����g\Ā�8��~��HAN������縄�4�2o{�L;`7��w�/�Ԁ� }m�T]wØf2�hc��l�NRV��
��Fv���;������mi�o��=�Ow���k�Ćo��j�f�9�N�����n�xl�v���j��[�E�0��z$-TY<�H��p�&�h���h�9µ�A������+�m�����3���φ�4����P&K��.�/%�0���rN�a��	�NhH���,i)���x*^�N�fO�9�����䛃C��$7 �Z����-[�F����\e�!J������r�7�M�C?*�凒�j�ff���sxG�I�9��G@带�[at7�X0��݊�,EL�����'Nc�U�b�'�ɔ�G�j��qaAk[ /�!#�\@Gd�F)L����%�3�$,�X�����ғ���jp�U�Ӵ����m�V=K�BfH�}��:�sg��亰:�[Vo��oE�1�!F#U.2�ַ�Y��?'�y�v�r��V���HT���OI�L#2�#��m������n� p����7K��FE'��v&�|?�un_�7�09�T����?��G�Q� �?ĝ���O`Q}�2�鄥��H�_Y"��4��ԕ ������t����/Y�mf��wVt�0%	J��lT��樂D�c�7`@���!�Z���>J {'�"�Z:���Y@�-�PH�.�/�Y��$t;������8���Bo���3��30�fu���H�Y{�+uv�-�VZH1&��L��콰��c�i����N���#㭱���J�AI3\� ���ϩ�uZ�E`˝w7�-��6�`w�������6�B9O@C�!��aQ0k��ׄ��7@���z&^4���Vؕ�v`��xܫ?��,��%(d�P�k6� ����lp���m�iO�9B�X���\��}#�抶d� �x`�W�d�9�%��a���	�h-p�U�߈bu�Vsq̛��e:��Q�q�����4�l�xc�B����ڻ�\���+g4�e��P���<���㥀"���;�]�SM�ڃ��]���yq�'�L�[��0�o2�֪������JW"��2y�KE*]n�ժ� 7G�!�2C����`��P&�>�����W%j!�n�^�̰%YR��x��֝:jݗ�Ι��6���$2�D�G�Â,J�5-� �rՍ{��Ɓ�^�g�S��L����{����uO��a�BXj^n�:j�0L��J����e:w�m)�C��
�+��_�:������� ���x�����m��LS�ݥ	Qz��J
b�B��y �kJnJ=^z�M�y�w�h?͎aq�4��YL� �W��ٞ�W������s�˴��ci-��z[	�O	��SaF$����SOS��c����O7'3+I�Q�%9�hѧ��4�@[�<�L�X��=6��Vi�9��ڳ�/�#��w�k�xZ�D�@1�]�̏0U$.�})���p�ou�c;7�K��mF��vՁ&AF�)q��	�*)V�M���2e�2�6��#V�?��^�g}G��b*����i�-�~8cC�Ŋa�����򎿸V�S������Z.=ý]S���:���ߴ��=�B�Z
�РQ�8K�F�F���_|��@�C K(�C<․h��^yi�_����������j�\]ձ X_��UCWR�g�acs�Z<B��
��i�}|%= �
�<r!f�Ui+.����r�c�/�-hk �-Nf˹@������ ]�'%d+�?&�7Z-�5[oW�q�?nt�ym~�Z����_tpȱ<�PF�*ɕ�V�����2��H�a͆f���d_7@����U˖��E'Ѷp�Brr��L&@C-��.ex�D�E��٪�*e��ta������[sǲ�BwL]��}��ՙa����U��`�O�	�͝���KlƂ/��E����'xV� ��VW"P�ɇ�7T�����'�JJhS>���_��0�I�m3���H�r�щ(�Y���.��V��܇��2a��N;�>9zx���������<l}9�c�]�YZX˙_�8�� ���PY�\��\U3�8�G8��ɟD��Jᕲ���.�ޏ�Z��1��b`7�Q���4�Mc,A�k�R	E���@�Gd�wf��a�=FU�ԅ��x&"l����{�	�ŶR�[�f�WI�>9��=z�v����d�|��1]u=b��A������GO�}6�VN�nAP����6$1��}��$���-ud�J�[��$���_?cO[�NA	�ݴ#���3�J��?Iu��~�L`8�]�\{*|uV��Yg�G!Q��] �xsy���Y��θV�b>���[
�~h�Hei����ܽL�&� ��=e"ѱ�ko��UTpEojD��P�%j�x4�B��w���4; ��W��A��4!1u�?\��f<g�am��0T4t�L���/�^��Ѐ�N#����g�?zH�+d�߲��g$j�m��ƘB�5�=O�x��l�C�
�I+�% �l"&�V<�s�� &H`v��c��/�5(k�C�Fxj2R�'�~[ �I�j٘��R�����"nZX�(j0��h�p�HP��C���N+n�O��D ���-����ZV���<��1H���L��qB�`�f�Ƥ�\��B׏s4ۗ}�����&u>��^ƭV?�$�se$$4�Y�ȑM����j]�G��ꐙX��%�]�k�z��t�35�L+�׊PZ��,��w��o��W-�Ȗ	E��#BY�l��\�">m�i���5��`ݖ��ќTu%W�Ǭ��+Weݚ7+�&-��|�ϕ��ҕ�L�5�mD7k����-P��O��b@��sw�o�+�e�R�*�]P���`�3T�ϣ�x4��v�M���M`��0�xA[G��}��s2 l2LZA�����o7���%c
TT��RB�;�����\����P�y�������ȘИ$/�����HK+l�݀Fw-��h�'�,*�+~�S>�E(8?�5vxl��$�uDjg���
+�˚����Zxeha{���nK�dO�X�d���#��y1�#X�X&k� �e	��<��%�]�@��$D&H�-&�떕�'Z˰<�T6[�I9n���Tߔ����pp$�MS�E�%\�82jpoQ�զ�K��-q������MI�t	q�kA\u&%�`6[��)epP��M����i	�P?�r0�D��.̪j�z� �u����L^��7Z���'�̲�I�]�]s�{Rxv�lI]Č��a�X)�@������T�f��
'*�z��������I�N��j1��NV[�1ր���m�w?S�`�7r��[�N^6�
��,9�j�����C4��*�'�_�%�r�y���|�F����c�����]�.0�Y�h\ݒCwr�[��vv�-��~z�ZN�>Q��K̜g�;�
���
���#��
7Z�Q�����p��C�J��A� ##�D����@r��6n�VU��`�5y��E \���)$Js���Q3ȡw�9�3o�����#p�-��BU��"��h�����Q�L���c����S�Ҟta��ejZ�0��i��ڹm��ud�t�Itc�q�S��1��j8�]ҵh�^+�k�@L�>��	����u<wUy0[W��%��	��H��ǐh�\V�/��)8$U��u2��3�����>�C����g��Q�t��x���p��Pl�J7�3�/&�.��sX)"��Ɩ�D�ؖ#3���tx�w�D�9���'�7�6#o ��Z~��½�Qaz���:�F�;�D ڶ9z���a)��37��A�o%q4O��u���1@�L��m���Rp��{j_P^�!1��?���s�����X��-}1������wF��!/��OSM�kda��_J{��+��.�&��	��ۣ�7��vE���˘��3"�u��tBM��>��M�ґ���(��aMPLs	�k]�A�;�|<��ȷhk$�*�LV�i��v��3�a%5Z�|-�j=�'7�q��׾]�K
�'�9�9z��
e����R ��1[��-��^9�SD>G#�����jW��]UgGs�����_�ʜ�"'���6�ә��� G�©��g������,CF8l*���|;I'���9v,���q������z���r��%�a*���A-���xLc����8�c��1�^S�w
l�	��r���������:�:���@9�fA�;�}:&W�N*@�J�O�(6�����H]��+�J�*4![def�	Y��3w��2�;H*N��Q�����W��#	|�7
_bcDw��{z�y��l]}��e{�U��͟��#�{���"0$���m<EIOw�vJҪ�		�!������2�biT�Qa yh//��*����I�g�ޏ��nP��tV�V��VUMf����~���
��%�4\d�2���t|5��3<���9�6c�;���)�ެ�C<,�ԫ��k�����)Su�1���m�Y����ę��L:zV�]#+�Q�t�P=i��T��n@��)�:?f�Z����	=? [h�)ǿ�h">uG�)��V����?ʧ*�6M1��䳈��"$��D�.Y3�"
��Re��/�?d�X��{�0�.a �'�(|���ٶj��;:C�O�H!|Ę$f��C96P��Z��4D�CK+s�?Δwx��ap�>Tu�k���U���@�a��u��U����lJl�$BF���ʆ��LQ�N\}c����J����f�ۺm�PLuCa�ۦ�����K�a���)���_����Eg�PxF�"�!�o[�jK;���b�-Dn����C�T��'j��_�2�R���a�%��XET�b�t2��C��t���к�i�?xk[��[��h�s=�[�~S�J�8���iX-C�8
�a���=��p� .[t�t��b�A$�눋��F���(Cό�j*[Q�$���37r+G5%ieX+;f�R��+i�0� {�d������0j�xЊ��ϻjӞ:l��L��+�ՉX��'���!��P�79n$��_��RU����W����+���-[q^H��=p=���]�8����ybr�3ǛR:,�`Gql>��SR22���=����-T�%Xf�S�'>�����lK~�{�j�����>(�f��k�\�[�S#��^A���.�i�L��	(7�7�x�s�A�����hcMUdR�}=T��-A�_������*}I�J��A�GX��xqkb
�攇I�v����Bq��7�ͱ�3�4��r=�����l��y���6�G��^�)	S:�
 ,ʔP��Q\e�xc����I2�yݧ�:=��ݠ�	 Đ�������l6����ǩ@��"�^��W��A H����3��m�6͈d�fY�i���4��=��1FF�iYz��-�ޞ�(�>O@���V��z�uD�V������H�Dq�6j�z�_qpGqCn�s�q��H�ƺcM8�h&p���3'�(���;\|��}���W��y��i}�9��!*�ႇ�(�=x����i]C1��FN��(d���S:��ۦ2�^^��xnj���hh����[g���ݲ���Ŷ�i��Fv1N�u�=��D�%�aJx�/r�O�O'��䪰�Y��RU���� K��&R�<�
{މ�L��m>�G�����P�#��"��̢w1�f2���L�h����Bm|"��x�E�������<�6�^�����P�Q�P��?AKz�q����Ec�'X�|�|p������b��ƫ8(���\��A�ֺ��Y)k��S������`�U���g�<�d�)o>�5���l�j�j6�0��ޮ�����g0�泄K�Ў��tg�Bj���HՕ
����G�y�)-�R����j6�+�EJ[iS[�lu+��d'��I��U��AWO�:���YHt��9n�\j��ZGA�c�~�Eo�q'���O�?J�~}���|�Z��w�tcZŝ�ԮPJ���Fu`b>�^�/u�T��S�Nˈ�� )I���cbJ�=�q�].��Yӎ��2|��f���lB�_oLI��TG��EߨP2x8�s�%5��u~��$J���3E�Y�<���PZ��>��$!��5n��$�!�&KMm/���FiA��"�S��$7]��LfP�{���N��A�z�{Rn�M�B�vC��=�[A��+F�A�Dbܼb�(O�ey�%Q��t�x��u[ ���� bJ$�@魧�4��ڹ�(���4!����
�)g�ٸ�Kq�㙱#�;~BR�L�P	fY��A/E����9��g�X��YZ�%��ް��:<(�w&3fn��_�M퐰�ݼ�d�^�D0Q-�f��U�tyagB�tn�zh��/3F�5q�#�z�B�����������G0>gƨ���~r���l�;_���{��&�44	�hCU\�m��������N�E5YxD8Fߴ�ڮƄ��'Gq���1��/��F_19����r���M��\�'۟PP�~و���tA�v4��P�`>��ްP�0�d�ݭ�Y��z�d���� �6��i���?��]��6�CZ��S�i�T�q�&�}9��ڤ42��1@�.j�Loe��j�h�u�买O$E��YN[���G�9��g\��R��A������o��X��o,�$��I,3v��aj��?�Ȃ�[}����Ļ� M�S(���(߿"&BMS�e���5|��dH$�F�j�������y̘?e���F��>���jT����G�J#{A<m�m�lU1�tv�6�����G�w���PPK�ֿ߬%���k_��[ �(�#��p"s,�wȖ���U:'�C��M�=��cvXO�dW�13�h`��5�G�I���T�k�ӷ�?�E�Kb�bp ��D�HQ�P.7+ƙ�h�r! {���O��w���Z�$�~WP��|*�to���N�?����o���GB,aIJ��G�]���Eْg��UX~���5�3/_2v���5LZ�,<M���Bo:k>��m�a_��@vO��u'�!����g��,�b&nG�/���o8�_�;��gV������@G��ۻ���V/��l`kW�>���O�}?��Vt9��7�Q:����F%�d��$5A&0p}?O&����t�o��y���;e�����.y>S0'�� ��o���[��}Ï��n���{,ȶL���z%�(�P��].{�� �T�b�:E
:Gr���>7Y��]ΖU̯E]����Dpђ�Ν�H��U��,O3������Z���i��5|�wWM�QUo���%��S��4)JgduM�0��p \Y�d	��8_uj�"9����x
�6�<	���&��u�QB��d���(n+ޘ+r�<�ʴJ��_!׺f��E����h�x�By��"��������'Y��ΚU�<,��P�}.���}k�C���iu#�5T`��(�w_Iu�ˏ���Z�:��B�d��̹"1m�=��O��r�"m�����X��^�Cw�	��e࿴��� ������*xA.V��3,!���,�BD��^�� ��#_�7����� &rIP�L���[�k1�n�eÝȚ�xC���r���<�t��HD���^��I�a�!۝
�	^Z��]�.Y�}�M��%q6��#�© Ͼ�E�%U*^�5��
��mV.@�J��b���B(���f�T���<]H*��=~B�+=��9-�X�|��h�M�/Mlfن���T��NTU� tE�oMN���7�L��9��W�D1;�]i[��҄p @���S*ٞjM�.V�,�ME��?���e�����^��m/�x#m��%T�D���F8)��]C�۶��έ��Δ͚۽���S�{�V�A�:x!͜�o��
-Yd�Dm�bVW���?`r!��n��]��|9�x����5�"���h.0�(G��☦���A;MTٰ��kb:zD��zܳ�V=�c��Y�X�˱!�9AbP�;�5?PS;&(	J�n�����*�8�[ ��+�$ܝ0F����z�I9��?A�k���u�[�:zհ��s��Zo�ƱT[���ǎl<�|�uQ�p�ks[�rq�=JS3��Q�}����NƧ]�.���ln��T-@�F�y�|Cf��虊t���܂
��.��B,9|��΋P~/)��̃xV�
�{�lk������%��e-�+r�MTA;�8�Pg5k{���5L^!I;�;�X���zF�Z�f��xg`dyYڒ�wO��*`�d��R?g����=v�SaA�?�j
�ro�v7(�����h�s��R�|��Y�-:h��V���=EB�53�Go���X�>�|h�'�'�6���|��77J��6/}���:��O����6�QA�.�z�H�.�^yf+Ւ�R�%�z��7I��������}���=�<���p V4	�z�U�[��t��c'�z'J�XC��[,ž@^1����x��1m��>Nk� t����[����[�J�k�ƈ������'9�����:=섳Y�����<+YV�8�p��Һ��|Fp��`�P���bz�-~ �[��iU�n���o��6�dU �i����%Kr�K�8T�t̥uX���1���T9��g��ALGa�i!�H6ߏ��bl����Y�r�`k|
k
�dd�V��ѿmB��ə
���R���l=#ӄE���l�6�Jp�����O���J*
5�|��sɰME�&��0�bvXJ�[��"�ߏr��Σ_�u�Ό�����+`B��L�}�Y/��;�	�j�_JKD�R6�i�F��I�r*�g�[I��ik	�[e ���֥�Z����<xP�b��:�pXeH|�Q`��8��
l�5>��
8I������38t@X
�Csw���@��"��2A��*�\�;��.5I���)�:���}-�G�����N�漯>�(��k�p�6:~��1R����J�PV(�� ��V��i K}�
�f�x9�Dպ�@��:C��1@q�;59�z3�\`��6\6��+�[�_u�W�@��$�V՛�j��_O�,ho-��V�g)�����-;�cFў7�g�k��>�I�� ��֥|�+K��������B>��V��._V<>���P����_�Sf/��	���b�����r��@��W�,��������"sy��p����h�~���,N��, ,�P���YHu��{C�@�|AG�0$��O���.L^a�+�2�&��e�Q2D��7���8��x8�T��c��3/6ȼz~6�13m���P9��?�cP�6C$;dp�%ڬ�I��-����,�xv������2������^�>֫����}��3@��+�J�F���0���8���Nko��C{7K�h�B��|���}o��9��eZ��u��{�#0����6}�hrh�>�8b1?��1.�b��.W��"-��c�O!z+��$�\#�i.\&HR?��A�85��K��j��V?��l� ;hx{U��Rt�����i�}��b��_��ɏ0G#B[��k�@4�|~��x�bic������xuD�Up�@����.�s� ~��k�/��^ȧ�䏣,�1ԛ��]�cx�E�Ԁ-��%�]}�E���Ey�͜�|��:0ĸn��}���pw��,��+T�iH?׊XU.���S���Q�h�l�"{��N2���,�F�CX����U�8 =%�)�ü�vm���)u�H��aCz9�fz�z��x]�� �.�pa�Bu��:P�e�/@��_��K8x���U�7�[){�	zACjM��Ϧ����`-6�����V��_d��n���k��`�φ���T��q[c�����݉H��y��_%�2�6b&h�l��g���Θ�X�us��_���d��&�f�Aѿ�a{��	����?<�O�m�h�����ig�E�	�!�H�! r�,����U��=�Ȇmt�R��gfKHm��߷���5��c�oʾ|�@�spt\L����:��p���Hp����8Tx�9�R���ե�Ï�+�rʧ[gp������ 3��<�	z�d��<~|7Q�Hc��x��Y3�Y�OQ%�)�@�̟�_���;��X��EPŬ ��3))9g�Ut�ģrލ�W�c�t�.���w�ښ���qo���rSM4��i�?2`W�/���+�1A��S�����)G�,@09C�(�R:�rp��{�����ɀ;x��^��R �[�9_�ϡ�:ΦTT~T�և���JHx�����SBz�j
�=P��W��� ä# Zǎb�G�+�3��Z��4��}�����k��Ȑ���F�
s
ܒ��f�_�s�̄�i�BPimގ�6���
V@��ٟ=2;���J�� ?��
�j����o�`�l�{�N<)W�b����R�K�����1�
�sl�������RC�H�e�{=���b�(6�#�Ǩ��	��p[�u�J��E@/�u�q%D�͢��Wީ�1[�7R�oG�*l�Y�f��5D����ҷ7�q�{K����3�^�+K5	�%]�.۩ p�6���-@?�Z��H�;�VG$�4I� `i,u\+�������Q����n���
w�g��=0YYSf`�IO����B!D9��8�/��O�h㌖�͠q\���m�F'p�*ש�6���̹�L����\�oS*������� q��D���P�B5���[��缬G��ܯ71䘴�l{��<~�Δ����k�մ�I��,4�66�%A&�K�le��[��Hd��&��i��4��\�8��kl�N���#��]����)�����)n�3��g�V�&�M�M�D@p�Gǽ�.���='2,���:�Ⱦ㿝����=�&�4����]���JU������������!.W��-롴�n4�.$�H � 4k���\�#�Պ��p�J/A8�;t�AOS���.Mt
��3Ȑ�+��tj���BsK