��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����0� ����遼�6������"���#�{A���'j�Qj} �}xT	g��F����a��f��洜K%g==�Z���L1������bG����XB�k6T��w+F��3r1#�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>c��mW���rJ(���/	���~J`2F�x���4W�0V�y��l]��X���8D�G$�ۻ��c��rk�E8o��W��z�����O�Q�F��?-_�䰹��Ny����o��:���l�,�:^�G���G��ta�`����k�G=O|�#�ʋ%�����vao�u�_�(���|�
�O�:��h���e�!���d{Ϣ���
�j���~c�'�Ӌ$�M��j�PAӄE7O��Ε-��N�������M��#�$z�ވ�U�
��iт2!_
.�c���EwKgP�䷴.�>Ly�d�-���/�y��<Ûk�O��=�Da�����_eV�B������7�G#�U��L8�-��=3d@��h��e���\-	1�Qu$�.;\���?��$n�E���^�w,�m�C���_L]ѧP�M����\Pk��s��Zҕ#�_5���L���-̫�#�nq�7-hd���t$3�u���sE��Z}+�x����o��j���}/�Q~����@C��)J�g
F"*�;����H�(��.��{�������,���91�oƙ�VG�5���G�3r��h7��t+H��>1��
�5�uD�c�mo�����i}�P,5�������``l%s"Lr�9X*��޿�� |�M���M8A/�s�C���3V����UVa9�`w��E�%k�s��:��fí��M�Y�G�A���dQ����L�����0̶��tR��+K���R~�̔��q*��>a_�}y�OF!�Q�kZ�x9'�mw|�P�7�L.~���K�7:j��p+����Qp�2��`n�m�>�� 57Sz���is��\P׵K+��-@l?*a���w�1ц�&X��׶�(���2��T��s+�[�0�0��Y�z�*u3u�������l����O�|"Qx�0=�OZ�"�
L�<�4��;θ�mwd�x:��<AjC��J�4��r�2��c���%�r%<�3j���z�c���L�:M /���D�VL�X� gt/����6h����s�3�u�0�sβv+�I�ϗ������+h�~�u�E�E|�_�R��\,{_bh.�B.��{)t��~7��^f�W���/x��^^!j�+q���v}o�#�Z��6�lkw�b��v�
���-i,��I�z�G2��D���l2�aRU��~�����aձ �)��Ί{m��O�����;(4��S�N��DP�?l�І�}2꛶?t�H���4 :;�}^-ij1![�F�Lz��Ҧ��Xɤ�}.˔��1�7����;�u.^�NBR|+}w7}��e�7dl���CV���Qc�V<쯲�����3����?o��^�8ؐK�@O���?�|��g�x��������k��ET�b�mMK�71�u�g����o}�Џ=۵]��E[�J.�$�<�b���؀������ ����'����V����}3�~t]���Ѳ
����󞷰y�LG��f��<U&a/���{�M+q=T�\μa�����# O��ݴ(���3�:I]���C,ׯ�隝�L�n����J���1�n�+u�2+�+�:"]�I�"FA�b��ɲ2��ߏ�<���mb���,��I3>Ȯ�x�܉y/��a5�D���x�7��b�[ʚG��0���勥ŏ;��X�e��\r���O;�I�V�tS���x`{����M�Z��xy'�KJC]���n����=�� D�x�O�z��j��bϰ�JM �R�jS -��D�c��.OQj3q�~��(8�J��e���=ecN�Lj��2�9ڲ|��ӑ�V����8�=�,���3f�?�97fxQ)E+_�Z����3��_.�q�a��#o���:m:p��~|��O��7i��]�y��OSǫ�E�������%�ø��i�1��9,Cٶ��g�t�0��|��о��z滪���s<��&'G 	��Zt��K;ྜ��I`�.��V��r�i]C����A�J���?؋XR����b?̑������t��Ke�����w9�ԆbaM1F�st@;-r��%�tU-�^_4�=���F�-�m`��C�^�g>�9�p27��D>���i�k�R+Z�:F�9ύ�d��4v���MY2�M/ ��L����0�v�Ѓ�q���o��Ĩl{�˴Wz�S��3o��=�s�C�L��2�����5�mEe&T0R&Ѩ�Z(�,�a�GgZ;��}"���s�Ř~=�G��^��'��_�JM^������t�Y�*Vb�z��)�B]P�Q�I���i�x<��8�!$���;��U���h"4ø-5Q?���o莅NRa����w#6�#"�%�n.]�c<�r��E;aS���(�Ɖ�#����)���Q�j#�Ǭ*.QD�!��e�������G~�3#ɀ�k��h㓶��`�͍k\�
V�݆q��'�6��R��t�Q��	�4���s�{-���_Ӳ��4�Wn7a��@ r��?�D�1�O=�^"'&�<m�?.��W vg�b�q)F�=�0j�y7[���
Y�5�pH��T�kɒ���G�GO�<���t�E�Onz�Yݙ��N�8"!��ye�2���b�ǧ���&cs9�A��%غ��]4�����i�ʶh\Ҿ��"�i�N:O7^��'kZ1��'C�M�F%Eݤ�|�%��,2���b�b���u8[]ZZ�{�W�C��UU�'ܜ�Y>��~] �����ѳ#�2���?%���,�Z?/��\�:>�HL4<$ޘ�9��1���	�
�v�&��㓏�W���K����7[S��[������j5����R���D����m�c�:�}	������#�����&a���fX���[�*$8���#�H�f�=����DQ9���MP�f����v�e��PQ���$�y��A0�U���%x���b����pG�(�6���j)�4Ҽh����)X'R%�����X���1���~ԺC������F��3}��K�K�_g�*��)>�Eҽ$����2AMuJ�n���?�@�J<�>38k��/�Wo�����V_�47Ua�g(`f�gJ�k.����*O�\H1�ײ� �>Y$�9#�̒x��)90)I��*a{q����1T(1>�~�7��e���-�2w�C�(z��}/R�� ��%}�O����LU�[�<��J�0�u���+��ɖCf�A�N`n����#��r���a�����qa/m��}�O}�X��r28�s~�q�]�-M�8<����E9����&���۲�R��� ���)�pL��0�W�f2�i�r�])0�|;:�g*���#:t���_���|�z}