��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���,���`�Q �����6�͍	),�6�md|_��n�x�"u������K �5owJh�E��qڑI9����%,%UEwf�x����;.�9��p3��,/�֤����"��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�A���0>�kz��/ �_M��<-�[a�%�����'(�S��jS_�,��8��T�.B߫C|��N�(ݝ_l0fS!��mYԥQ��DF�S;���h/��9mϓo��ޗ��L�%���QJ�8Ȍ��&i����_7�0����ѫ���'�53s^!c��׿�0���w�/aHc�^����b|�������"c��h	�,�a����#t��7x�oV�d��T�����|ߢ8*���P0�u׊���6|!	Ї��n�p7��t,��E�cV�o�����g�꠱�� �aݍ�����}
 R0��N5�b'�vs@��m&�T��g�WG\J.�{|�5��5�����V��#�ҹ�BB��weDL�4�p��~�6{=E"��g������_*��q�XƄ9����)�;;n�] ��׎9�Lϗ��Bo�T�@px�WQC�Z�H��`F�MWPuݯ0�ٜ����	�m����'���R,=+�d(@U��9o|���ۅɓkظ����;͎#�Kĉ��i����Ei�k���9��;X�2�Ģ���7×�ބ����R2.������g���Jh|� ����_�����������S�����<���2�P2�Ù/x�y�k�e�m��T�!��!�j��*m:e�͈*J���&�ED��n�S�l��Z�7���m�����dr�w�K�<{[�Zۉ%�&�i�����~=�ؠ9���C#�ꂽU��[k�?�%�C��O�����6)mW�r�~����I&P��n�����\Z!��V��ft?�Sv�E{�S��jq�%P�]�jer����c��B��:_��d��Y	z}#�z F�g��.�]�{}�^|t>��d�A���&3�k
a.�-@��-3�؉�Vh��ӟQ�r篁�p��s�a����llT�4OD�ȴկ�؜;�p��X�NL�R�����^Ę��7^�s��
eE8��нi�J�`�Эj�	�Vx0y��,��d+��0$nc��q���=��k$4��Z�]?�3Q��\.y�1?��_���?��{7��7{	Z@�+��%t��p>^�ͮ[_@_)���i(d�L'B�in�&i���>.���t���~��*c����*���+�#��b��ݸ���]�����AW0���>�����♔���O#��t���nZK�jA�2E�Vvx&1��� ��>�n�1�O75b�#�_���O�t]�jQ��^�M*~
%�Xx/f%�w"Hω�琓$��|�i��Vd4z"��1��Q#�9-D�vɋ��Q���h��·�qP�A�y(�-�����i���-�v5��bk�Am��3�D��1�1;9�7���jڥ���]ݓ�P�UA?�r������zc�Hn}�f�'n`$qV�,{��dAU�z�H��P�����YȿnS ��/�C̗��ݰLL���:;��&.�eɨl�Ul�o?�Qz���yU�@�^�ol;+nfG^�9B���]v)&*0d%�H1�`%5%�e'�a��ݩXQ@�\�w�B>�'��&/K�W"Bq�l�~��=�[��OP\u�RV��!�0�h����|^���݌+��L��g�u�9i1X�݌�I�ք�ǜ�86l��x�$�αͮ�`����+	��v�[��@�����bkHc]���<E,"���:��������m�P��O� �p�_|�Gh�W+��e]�����������x�h�
㴤��w�DF,���a���6����4��0�LJ(h��t_#���ζ_ ZZ��l�/�ɋ<����]�a��ŕ�1B"�ΣV��Ɯ�i�Ñ�}]�o��}��	�#c�R�MJ���a_m:���Ȑ����\����Dj����SFBt�g'G4鮤wSEL�|W�����HT��T��BMsܽ)v[�睥�AB��P+c��O��n���@�.�xLƄcu�
�}s�bx����U_�a�6Cg�¡�P^��.ʤ6u�m�u�'�!����@��#��X+��它Y,cs�>2�z��~	7:�JŵD��2��h���Z=����-�F+�`w*I�+�l�8s��ߥ늣!�2nf���;��ƛ�8� 0?6o�|"\�'���{X,ې��|-�Η5�=Y~�^ٮZ��K���P~z����Q��{�д�qw�1굶n���M4}�B�G3�N4����f�g�� �C���ri�\8g�3��?���_;T<�<`]k�K��G�ݼ��"�86�."�����lW;�&e���;"Tu�8�p�%�}J�]o7���(x�&�m�������E	�S�	��:����
;0�GQ�f����%Nd�yR��(3-v����7K>f7/ @k��ލ�l�Vu!����aܠJ�;4��?J6�$v����8W���xM��E����=	4ÿ0��7�X���UB�>�MaAm7���)�J��A���ew����ft�-r�t:?@�s�$���"#Y��ZЌN(�`�=���)o:;}�+��$��g��"��r�F�3O8Y��m�67�m�D�DCN��4����m�t��z��U��z��o�]�)���߷�D�Q-�.��1�n9��P�fє�����>�5��$)��P7z��c`5+9�����H�57��ź�fƑ�aCL�LƝ�a��4G�1Dh�o��)�ݿ�z����P�o�a�<DY����ւ��&�?W�Ny�	����H۶��	��lĹ
\�r�kQ�nݯ��k��g�R�5Z���%8�U�Ko�w����m����6��c%t�~M�ڊ0��e�O�Q��X��Z�	m7���btRe8��c�����y��ޔ.��գ���g�L���i2y7���d�H$��}���v��f�bَ�S�Iw���МԺ����O��t.�̺;2(S�R�Q��4�Qu+!�Ɇ����<я;#� ;q7�_�MV�S��Q��"(��
�T�b�p�-��X������H($�*-Ųn��U-���i�icq��_��w�'��b���W�2���*��S�	6v�BHjA����$�G����c�1��,�f��\BW�Rmpſ���;�����@�����֬0�N������lʉ�N�	��_pQ�X?�wg��;Ew퀷@�&���" �\	b��>�^��ů�xv��� {������E���+�:�L��=�
V�,�K�N��[vj�QzT��^�iTZXF��d�X�F)�i��2����֭(|�#j~%F�V`���6��k�A����h@�|RG�"+�V9�ץ�ndN��s���������Iڈ|��k��yS�:�̃��x�p��H;�n���{�h�.+傑�F��H�,��T��6�=<O�]���C��=��K�s��
3�vW`_�ʨ��0=����#�i���z��#u��8m=�wC8�;\A�O�u����(������zG>z	(�Ȳu��ۋ���Xn8��~��7jhQ�`��̖y�0gB���m�}����{@f�����x�TS����ok�+�ޘ�z��X)rg�8U�,-J����aP&����ޒ���x�s�`����I�B�V��r�.T�I������0-���㝿�7r�����A�)�������y�Z���)pd5�9j}���ӳ���f�w6TD�� �!�q�.TyZ�F��[�9�z&��$d��ES��:ݲ"���҄'=�}�~%S�f3��!���%G�v��1��\!
t��&T�e��e��$�P�I��vcZ�^yE$��0Wu�X���4�A:���X�K5KO%�!�dAm�<#G�A;��\��@��_�kѮ��o��;.@&A�G�?�E�$��d1�ƇM8��+s��BN%�� `�2k�t�%��L9��<ؘ�t�D�Htad�� �Z����q���V����|��5N���,�2�j�ٜ�|h�,p����*(ݷ�l�v�]WM^�l�3�	Dѭ!H8Ut���c�sR�˵0;�0e7�1,��F��6/ '?}�g�\��W����+�9��Q�e|&p�هzG��� r����W��֯���؇�~ǃ��kO���vK0%.��=%[�mqzk�[por���Ohl�"�g���;�Я��<W���Qf��:�k/�P��^w߈S
R{�b�U���hp��(�"2�1v`pҍ��-�:Qx-�O�1?I��Y��1�<<�A��u���Q�V�0o��͏���Z�������*.	�4��hw�j{{�Q'D�?e��1a�����&�p�S��z
}�&�*�w@�څ��Fi"�n�b�O�-��цI
�X?n.��b!�u��ܝT���� "o�����iF�W�M�����^�J�N����2%�T�<,-�fYqK0����I�^�ċ Xg�uJ���<.5�i��pn�5Fq�csI��K���`!'Wo�����5-���R� ��*u�W�P����	���kʏ���K�c����	���@� :Ƨ����oQW��a�Ǉ�2��:�&�4�"��=Y�$
Qt�ئ�\js�-c�"��!ӻ��X�*.�Z!�ķ2�T��d�~/h�Y���BX�sQk/G��b�&�5b�uD���I ����񁼙j~!����RU�@tz����@�}Jɒ��F���e��8�B��j��pf!�z�I�N#�d� � I;���f�?���UJ��I���r�*W�V��Z���}�Nn�g�Go��3�E����J�K�O���]������ ط�J�f�{副������}��4���q K�'���[$)���""��G1���S���I��#�o\O��,�6BZZ���|���I6G+z"�Me�!}O�zéP�7<��t61��3)W$�&�K��n5�&��@�t��<��R��xL{EH�V<�O��<O��l�M��:
"9��Sz��%& �Rm��p��x�ou�@����$8�ݪ�/���v��,��&v�3Ъ��׿�}�J#�c4뤇��Ϝ�<�YnW�$�2��3����yw��^p�xU�-j7�����*���OCJç}�O���$.%�����XV5܏�n�O�i7ޔ��b��)�������z�|0���+�6��k��9�[�N��=Ⱦ���n�}2S��F���(��Ļ&� �X�8�m2S3��zϪI$h��.�V�9PY���0��C��5�d@���F.����Dr�q˸����������;^"U��6�}`20�Vxr�O���@'��bɤ�h��ɶ
x�o4t����z�x�v��^H_����� ��I��w��J�n��e�uq����	�[XHB�=Y�LnKso�U�7g��ǪK�Ç������i��ʜa%�=\�hP�t�[�&	�R\*��;gT���'�I�N���:J�H �����{""7%/�ζ�O �1rG��^����>�*W��8gB�ff��������\v|CSC���_���hd::8� �K�)o�/	F�l"�]���K�rE�����y���o�.����7r�.^�6�"N��ْ+E'[4�|��rM�i��F����2Dj�NxN��|Y���H����������s�6�4"���i�`����nm��V��pT�rL�c�f��a4n�s��1ް���J����J���_�̈́�WBvfQ� ��Z	sQE������J(ޮU�7��9�e�E#I��xx�*af$E>�쮸�+F����G�A>�)?!�Słp����_�ri#�R��9�.X��,kơ�d8n!,R��pO<��[�^& ���_#�ﴐ��;��.�n��7;���c3� ��L�^!�"/�l�/�3���#��}���W���H;�;�i2*��)����-�8�����[�F	y���^N������#�hZ�/[C[��F�k����OD�s���I�G�[����~�ga��Z,#��	�9�,wH����'���xj��NYB��-c/�p5�ѱ+���5%}�ptM��_�z���I����4|�a�o|%�Z���]���dZ����v��V��<t���1�o@Z��?w���v�xG�j�+~��b؞.nu�8�\ps�,�Ӽ���ư)W/�jǼuvug��`��( ��b�����r�w;��2
Q`�]��탍A+-���(�N5���Y#Ł�Y�K�e�#*�3�z$���1��������U��8�(+˺��|P�x���à=^�OQ̬�������6�;>�n.�/g���Iu�#�'U�HǿX�)�+�bd����~��)i�RRϒ_��(�=����$�Y��%+��cU�:�c���oJ����ύ��W�y�F��H.�To�r?J	BJ|���Ɖ����뉐m&_5����3���#�[(�ۤ�mq��WC�:�*3��A
�e-\d���}���#�l��uV {�H?��쏮x�/x}r����S�F��/@4
U� `��{���`498����2���Ux�!Cg���ki�T��%a&%+���k���_a6��[`�C��l�x���ՌX�(�>��l�R]�@$���y��Y(��9�GUu��r�{4���=�%,�����G1�����F�^:�?$�����j`���?�vt���}���SV�a�y9^f���UVT^`J��wG�R,o]M(��Pd�>M�Vq��@W��ʈ#�X���l�&���E�p��B�����G�h�����=N~�ԴIV/��h����8�rC??��O��N����'�:[a��M�9��0<�U��f�}�/��1�)Uz����O_�[ԃ���5�׼��(u�<.EˮAo���c���ww���r��� � �6bǝ��p5��i�P^�Y���i?v���m-�+�)�ܬ�L9��_��8E*�%�C|;kI���kX*�c��#��R�ئ��|��7���' |�5�K����5t�Q)ԙ0����K?����)IM��~�ȾBlzt�UB��6᠓Y�Ȱ5o����>'�I������t
VcFk��34�  ��s��C%� AAָ�[GN���!�r����瑝�Q@�tP[� �n����:�[0� tn+T氖�C]���Pғ�&m��������2a�:������;����SmC�?�RP�k�7�*�X=��]t]L������$����yw3��a�P8EDc.��='<�z�$��̺�J�T4�@jm_#����F��/?#C�bq���t�$�`<�2��8T����!����ò@:t����J��
�<�*?�� ��p�.�@? ��C�2�W][�׸�QF5�x��f����e��[��gӖ��=	��\�6�=�X�a��Zg�b���x�A!)Z��1*����5�v�H��<�E�������.��N6_[K�㝔d����-��7A,����އ�o~9�a>��1r�9P�I��l55�#�f�Z.�w+��T�V���2��?6�����E�3�O��F�<��'��%5�K�WW��Tocɤ��W���V_;K��۔��:>��-�N�����񉴙1�l��2�*�h��O�,ҿ�L([�5X; w3�CXo�����T1>���N~�
$��[�~����W��8�f�|��6UzU`�Չ��E�B��G�|�`�v�EE�!!�����  Ku?��md �{�V����Ҏ�i���ٌ"��^��8��K��@#+.ִq��"l9%Wc�cwƖ:i��M�A��-�����){����I��iFY���i}�+{f$aD�W�\�)��/BF(��-��]@oo-�U�֔��[����BS�\1,"�5����i�W��T�1R��*}�C�+�$�M���	1�+9Vm��Ib���'��@w�����]�q�7Z���U�������Bz�o�Y)�����h.��tb��x\1�#�d�����$���`�%_�?hk��������/�f��,���ۊP~���9���^K���4`e��Ȟ�l.\�Lc�r[O��gV�
�k��	���������{jE�[��q?u���|����>z�#e������,�^�L)��"͌�ϧ�XZUv���M���rU%�6�<;��@��b�i��S��k������v#��<I騷� ���Uf&>~��{��~��w��稿��)�q�%�R�~cQ���fk��ͥ<W':���ÕC�Y�#�m�^�]+�χ�^��0V.����}��U���9���s��?�&j9�8�'�Xi�Ҍ�-�D\���/>����~�:���R/��G&5�4��q�n�O�j1�1軤���bY�*��z�	�h����b��i��d�%6�N>���q�[a�W�Ð��\s��PC�7v�ZVc�Cy"��/c�&zKo�}#�{��,��e�H["	�qV��͆���p��U�����9��m44�/���E�p-:�fA�^��h����;G𳎇�G�(������;���6rNT+=�Giե���I�|6p �x�6�J�e������� ��C��d�T$�$��J1��(Ihd��=$R��,3:�$�ФP/nsL�9l�_&����Y�&n��`7�kb"J]���-MJ���u#��t�����Uq�Q�R9O�ET��V�&�V����E��`�5�x�7���ܽk�h}�	C��\���_a�s��3r�̰���y�^rC;-8���hs��N��F<�j���%ڼF�rJOOT�\@�?7�������<��
�Ԛ��$��R?�J�cd�F>�t�N�ݳP���-���5��Y�8�	]��x�Śÿ���g�:�<��_c��nn��;���u���-��MVIe���1WX�g�^��(G�e�f�"�[�`���s�I@��j�} a¸���0�
�G�7QUކ�h=S[Fn�Ù���Ӆ��Р[; $.�x!��Q�o�Bo²wXt#��[W&�%K���\���D���L���O��	�|mȏj_;�����>o��e�z��x�My�v�w1%q:���x�h;���͐ʒ)���t����q��G���Os�h����fTC�{�a��޴����Q��{O�l#����eʓ[�4�Y��K�!~=�.,�C�14������eo��֝c���eX7GJ��f2��D���2%�q��'�F�u�.3��V|x>V�MbCs؎�e��	�N���St}`^��pҚ���R,&���[���5ia�+�P
^��?�{������C��t���mAfm�?������U�/գ)�̣�#�%��>��_+,�L�I�[ץ�O��hA��⼛]����D�:P�rC$���Nf�f���4�5�q�K�S4�~q�?��N�8{����K�r%��;����ԗ�\�d�f&��P�~'*����0��(�>�iL��g^�5��ʲ�����zu��Fטf��#u��l�0.�=���h�*��O�SO���s�~6�L=�d��g�M����)ƫI�v	,0�:�"�����h��Na���H���a��D���tӑ|��d��Q+bt�Ez_�8�d�����dH��/N"UD�эQ�7a�x������?_����}���b=x��O&��(D�bF�9��J���{ʏ�����/�-~:���L�C��7�>/��i�R*nEq�2+7�	.hZ�2��7�*~�����{�k��Y˕�=��t��H�Y��� �s�!mwn��F饎���*�Q;H�ڴ�J�t�fq  �/EKb�B¤N�vEz��k�
�D�^��Z��E>"�i���xv4'(Tn��܄AI�dyh3��%Tˇ�.�}Ѷb�s����Z��w��IE���s�^� #u����N�S�hE~�J$7����xq�y_{+j��q�M�(��@'&!��^9�b��CX�F]��,�i#,�c_j���3����j��PK��B�L"CB;W[�J���q1BRGu�uE�M<�"�?�q^���kn�`�\(������x��L��4�L|D�Q9ސF�a��D<h�Dn����>n`~�y��W��i��غ�Z�t�E�̋%׷+!f�р)�s^UNQp=mmӞ��U��3f$�t��5楟�\�P؍o��[Ʃ�ln	M�S	]�HK?o3:�p�ĩO	��ȟ�<��
ɰ���ǧ���[��t����Su����ż7�;�ӯ�U���{Y,:7j���8��x�$45^Lf�0ơq\�j������ʗ��e��M�{}��2��Me.>��\UHx�X|�M��X�u?����Y�ٟ�n�W3���Ξ�>���{A��
��s�;aȤ�H:O^�8$du�~=�aN�A�h��涫�I�	�(M�F����)����Mw�����HlRj���L����H=����/�^�^%�9r�=���q65�����w�/{�#�̀��-B0cMG�Xo����5�aNw:hj��r3�lޕ��j%QO3�_Y���$�a�o�s'�����Y�߶��Y��� �M~�|��� eBV�V�<$ZϽ���7#0���ma���>�L�Ju��o��ᧆ�tŀ%�ܷ�z_�|���5�4��=��B�I<-�Й�zbO$4 /⌹���a[�4Vp`��&���ʢ�X��?�h��;�#�_�ycΣ8��\/��	��o��Ǧ�rlIbBM9�?~����O9������X�z��j|z��8�4�C�O)�'������*�B�=�δ[e� wÊp���9g8�? ��F�����@!��X9�G����k�d�~l�V����?1���}oQ*�7#c|��okKH���\��D�_�����EI�����_��yQ�x����8)o��w��r�k�ϵ X�P�4@`���>�xd��Y'�