��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���,���`�Q �����6�͍	),�6�md|_��n�x�"u������K �5owJh�E��qڑI9����%,%UEwf�x����;.�9��p3��,/�֤����"��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
N�m�H2
��j�Y�?	l�Aō4�8�����>|�f[؁���
Ζ{�����0>��������'l�d�b�%#T���QOo�Rh��&42`�-�R3Ml]�Gq�]O��ל��J���('���Q�5�.����p��� 6�	J�/FM��8���b�)f�ĐI];�^�EL���j�����D�1�5�1�K%M6P�]���*"&	а��u��~ٷn$5h����k��O��L���׎D�y6"�  UD㍺���"O��ܣ2^ �4"�.��d_y&����V���k���ƭo����`���%ȯ��e��εA;�3Yй3V��l%U}��N��������aUiJ��������X(7:�_0�Ah9�[��=�2�5�����,�_���i+���C�m���K-?�qi�b<�-�a�!?@�3��w"�[^�J�������+��A��W�P���
�sYy�ŏ7j�S�����h����nK�L����E��#��-�\�9Ú��U���-|{s֒Ѩ�y0z�]�C �_@Jn b�K� ��A��a/�F�B�!�Ma��Y'�����G������]�LQ���|��gE���,\6���Պ�E?��d��򄻙���R88���Z�c��5���G��{,]n�M��������ܵ�l�{h�W�2;��+p�εn���>"q��N�G�T�����o�-�m�%�xG
�o�]n���	l��'��a��qB�d\|���Yc�Z�t�x�塳Lr��X��/'>]��59֥�'�w�ƣ����2I~ٺ}���Mw�q�ckg�<�B��<�� �b��ű�G̹�[�(�R����Dz��#hu ;��9�`6.z\��".����X*Q�dP�So�4�K��z�~�n�^�a��W��3	# ����k%��t��S0��9����N� �o�����.�Nj�z쵱�G8b�1?�v~�W��e�POOs!iъPU1��� ݀���e7��o��^�]F=c�59�s�+7�ҫv�J7=���z
��_�σ��y�\���h�_��s|��Z.����*ô�XE�@�L��:���e�P��E�U��2���Ἒj��iu�*�9*���^�y�Y��ja�3����qL%Q~����P�l8���Y����3p�V_�X��U��2�p�R�
J��p�ӥ�-�؞7�;���
����ԃC�B`)��Ђ��#�L.��FbOx�4��w�6�c��Y���ia�W�le�\�L����
NBR��@9��+����dϜBF�5��q�>��&�.{a��n��k��/|�i?ڜ��J���|�pP36���ҕޥ+�ϻC=�;7_!�g}u_�]�(��1Y׵��B��r����Z���aqB�������_��2����<�g�$��mִ�Ga��)�f�"��{(�3w>�R�5��D���t��8���A�����VkQl�"3����}�� ������z�����T�Q��@f,�V	�
�ib3-m�''�)5�4D���{�c�+&'��'�}9�5P�g8�����-;iaJl�$��W� Cǳo��zH��%N=����Iq�>n�0��| �H0�,�X�RhKM�Xۇ��tQl����Ge��j*��x�G��K.�"�b��.�o�\�����Kg+T�Z�����m�Ĺɤ�
��ó��&��)5�&�+�m,5TPY�Vw�~%8A|��=�H`(���JآD�ދ�(�K{B��ҝC:�%X�?� #�4K�������lTH�C˴�t�ԕ�(�<tۋ�$�� �?�R�o������|����O܏0qt������4����/a�+&[.b&����	�Vo�-�0�,�ɽU��-A&4�#[��u�d������y�e*��]�E�����1rGz�D�b���������?��C`�� �̲�	�Į�j�>|e@�T9�K�q-�C���7���C�kcn��DqZ����!d��su&������*��q5Ji�6�A�+�Ak�ŗ��Z�h_��f	}�G�@����Ԟ�������f
��kRN�������pm�bGCA:T������Z��ޗ9�Kl�
�f�ⴷ�����s�`�@����X4( ^v�UWP;���;75�U�
�\g�vC�HDM�&����H�i'�������>�M����n2fч$42>레Xɲ{�7�86޽��/
F�eQ.�~��O�rꢓg���@���!���@�:m?-T�{/����=�y7j!��#)_��A,gS{�G��,�1qo5աfK�b���БOJy4��&���\�Mǂ�zH��l>�`�J�.*�@SA��-��p���>��]ήq��,@�5vzV�����751����3���]��o��ڇ�P��D�d��l��t�3I"X�u,N"Z3���ҽ��N�¦g#I�EAR�>�!�O�cl{:�Р�Wtx��5�$�9���&Ha��(�F�ajk�#�:���c�,��f�A��,m�6�F�]%ү��M.0�%[Q~��A@y1=�����3p?��:
ʆS>W�wC>�vD�J`o�h�������|20t�˥����8G�{m+���m����R�M�:�葋�W� �E4�c�>���K���nHY���'��?Vщ�"p/�ysm�;7���l��
���&�W\T���y�E��w�S�>#��G�R�A�)i����5��CsP�0/�)��M�ּBO�D+]MW~V<��h�7/qZ^DqB���_��?��t�5��;��G���:�y����9)����������!b��ّ~]r"�j6���aA6�T�����R�8.����O)�Ļ��0���-TE��I�l��T�<��Ʀ(�G�&��	��L"�R�J�1���S��<�YrZ�K�q�l8�8TJ�e}�EbLZ�?M�[���j����92�rd�͏�n��z&Br��mV3���g��=��@�𦈇$^_'�8��e!4�g*��Z��8�5�KܢYJ�o����&��+[\=n���g��1u�0��=�1M͓FC�R�qz9Ƣ�)��i5诵���}|���C�J��CTWl#kFM��潋te�
_Y��!U%����Ğ�go�J�1�ңx�o��&jĽx!�������ɮ;f�:�M�tFF�I�?�\˜'�ɥɠ����;��ᶉ\9:�9��&U�y�W<�7���g�}}u����y�[h=b�-Tɍ�ND��kVg�7�@Jm��
�lk��C�4�8ÛVntY���yk���i� �)w�Ó����2��t�%Յ@��s�B/�/��G(��(I/�C� /���D$��o�S���
'�Oy��,*Hy{��і?�;,��h�����ͤ�O�z$��yqa;��}�|]��4*��X?#�]�%��o'��e�F�f����}��� �˞���N�G��{vOdf"Qe��w%��,�-�"t���-�e��9ä��wa-c�Sy2JQ�
�:e�n����Rx�#���qڧ��\��?Q4^��W��QZVq߭�O�G�?ᨨ��DAhcA��|j����^�:��X�B��(JY���Wn�-y/L���k��)������ϥE���~����`���T"�FJ9� c��1
�pI0!�.�|ZXeޔ �"� ��.!�m`�Q�Y�{Ri�?��h&��ǁm�Iզj�ˮ�uUlB?}w�j�����!�����R~�V��O(�v0�F�����	�R���ޅ���Wd��N�G��
 ��Mn��"�mȿU�������>��l/ӶSg�l���#�4��>}`1�I�F���V��;�iC�n���j�~Z�A�&�]���^ʫUݜ-��AlOӕ�6�32f�wo�f ���H���i�o	ߌ��*�U9��q|-Ɏ-�(�p�/˦2"���ࣦ�c6UyB�n/!`�^�_~��	[��D^�����3�@����u��{|ux6��KÍt�;��
}�w) $�������hY@ m_�]����^-���	�q���3����oy�m�)���A���GJ)��?Mo�u<&@֝F�+���#���6��O$���M%����<
P���̖ѭ˅E����O;h�4��VM�a5�"�=ts�2��*�g�=�;�K�je�̝���0��Z��:e2Z�� %�D�I�7�*R��k��!i��ϰ�Ԑ���C�6�J���cGŁ`3�\h�0z>���ˬ��2��t\��:<omfǥy��|�}V����`�;<+_Cc�ʁ�,ǆkE��{��d(�q�+T�݀2^{9�����m����_Q*5���{��1
 ӻ��^�:_��{&�U����:����#r�U�"^�*�Έg�[�c����C�$��&���4<��dD�G!?!���K�At���_'�:�t�R���V; Sd���1�SQS���>�&3�cJ��9�����[兎�a*KU;f��i`�3�
C�]�Z��_@*�\�$�ْ�v��J�r��@4ל-�p��0���]i�RH�6Au���R��(�j�V^9�)��3^'/��)�>�na�c���/?�U�\OaQ���U1�ܻڤ{�	~�x�b��R���+8Ҭ��^���qx�d���Qړ���Q��Z�n,�2�8�mS������)-)p�a�
�EY�� �֪�2���X��7�>\0Sr�����l�~st������ǯ�3Ҫ�@�:�����6�c��=����MO��?س�sZU% �y���1̉�}�E����\��cZ����dg*"��A�2��
�(1ː�\u���)DԷ���s��;?A����_E���� v�(Q6� ���LM��
�O^
�ͱ�4�I��`� �D�T�$%�Q�]���F]I?B힟�-Rj�J�Yɂ?h�@���¼z~-��&(�/O�>�ٔS�$ˈ��H�����Sw�c�P�f�N���/�ڠ��x2���_�;���c��b
 ==1�tܘ#-�*��6bθ�Z�4K��O��Һ@"�8ѧ�_u.���(y������ �5 ��p_�.���-9-�׹v�fn.C�F�fZ��Q�S�[��<�"�X5o�^j��Hmv�G{�֡��8�E;��1��`���{��]�����Ԋ g��z6J�3��
m%�uh[T7�%s���$Ķn�os��k�+���kS�p�j	��#���u�s1'��gU'�1G�3���o���V�ֻh=KkWK������lE��aDU��:�n2�y�*�/Hj"��6��DG6+�x�=Z��B�0/R����AVz���xs����)N\ε�w�8�/�ۗB�ޕ�/�*���V{I���E���Bw�����4��6Ri���"\ɸD�eOr�8j��o�W|�r٣mr��Z�]��D$ǉ=�p�	�Z�n�X�:TɍAG���9**ܱ����b�=r�
m�S�:I��@c����ڥ���A|�e�a�N$����7�ms�����8����`�f���$��-FRJޚ���f������~4$yШOkO��e�ևx��b}� *(؀"c��XXQ�J�Q���?�Ņ��+�^��mt��0[CV������wt�X�g?�%�T�Ѥ�e� �y�ۏMk<�U��m]�������"�E����@�lr��'��x�8�p�z5 =�,�7�?L��f�(�l9X��rG�є��%,�G���' �.:�����_1�@ڳ6�����E��`�F�3LJY�Xe �ۜJY9���zEjd~��^��MSn�^P4�Y���ȸ>��#��3K<�*���y���G	�?�}N�z*26PG�ٻ��,���1���wdgu��3��E3G�{�L����uw�T�~.Pv�DM��QU��,h��S`q�c�t�ZGX��'��M�ӂ3�m65wH�$PZZͨ�_,�yb_j-��@4TFG%����x�h�!��]0��ؕ6��}�^r��~W9Z*�V�����q�/Ո���4+bP�����M����*%u4QDϸ��M�4p�oB��t��6�#W^$' �O������4{�%aY�̇7�u���K��^���ms�p���k�\��@�J.6��A^��_��Ϻ�ִ����5�=�
�3�{�NxuN�!�޼��Yj��Sj0	�#���� ���Y�l�en�pN�@�t�(�J����%��YM\�����Q`=$�י��@������|�I�dC!��( %RY\�K��)?�gd�2y®L��W�<���MJ4
����ĕ�T��Lh.Ţ��X[FrK&RE[�-\[nO�h��c%�إK�����'&|W�萅�F+k��"�e�J�2���5n�:�˔�\h|�]ڛEU�{4'Y��qE_*nvh!���I�g�̯݇�/�w/v{WFH��R�8��D�U�_��ϸ��d���,��&��{�5>;��J�������xG�*,�s��O�&1�>U��$���yT��W�����A��zC���*L���1�O�4(���#�f�S��Ў[Z�䕤�p&�\<�g
�?dZv*�$Ye�W7i"���Fɷ:,i�]Yl3��T"��rYͫ��'�pp�y���,|i�i�y�<V���3��ٞV�Oy���W8.k<����׸�Ʀ1CI]�&Eb-��e��N�+������C�,`��	��6#�xY�n>jG��(�^����+�S{n�nb�A�y����Q��9�e���+�APv�ߪ{�B��Z����e�l�P����=��B
w�:�!�X[�ۖ�:�#���@�:V1k���$��`?��\�0ə������+4Y�[�����0�Ÿ�m�KI�4���6Vj���Z<ͯ�Q��E �7DL7�?���44�Č�8l�%X�D�"���:�J�ѬǸ�a��l$!t�	�@=|G/>J��-Ĥ�Q_~��6�U��%b;����3 F~`�Ņk���̓�a��"qV)Ʋ��F)ڣ���
��<�UĐB�)5�l7qT�������g��O�2g�>+��O��z�(�[���4*�%��kt���*�d���~	@u���x�M�_�fI0>�d o���-�oa�e]Pd���cQ	̎���Q�9�����G�^�~켷_�j �.Y�-�[�����O�r�����&��j��{�����s���T��)-������#�Rf���*�;\�w�[uY]g����I�7R9���fཌྷ��#�x�S9�حޥc��$YΜ_�n-J���=:����<z�cYbf�G�B)��^.��� Y�_C;J����
g��||�� ���W%V�5��G���F�f4&��i����հt&'��H�2�ዥ._6%]1@�v��
��x�RPc��ןu�<�Fp���k!4���{Xl��ӯh�Ӝ7�n&v�uJ���!��qa=�BΊ0^����	D��v@�׊2|zq���ڜmq(� Щ�%�A��O3fYgb�Y0�*��-�/��t�[Q��(�1�4ટ/���,tu�џkhj��5s����ǥ���Q�������?�ˢ0������F2/1c��N���[$�j�9�Rs.�l�j��!K�B�S<j�l��1/1�z���>Y�~��?x�Ѕ�>��U��Wm����Ob��S�����n�4I��"ԔI�
� ���E�G��ڪk���Uh��T}K�[9�s[bA�t
MԮ�󏡂��A��Xd�G�Ny~!Q���Z�Z�ś�2�u��JQ`����!��xACi�ڰ-��?��TV����+a�M�ie��ui�p��k�M��0�f;퓍|=�- �HC%봊��a�w'�;���т�	iwb�c��I�[�۹����c�k�耵��VCx��:��x�gs�uV�=����/���sJ=
{a�a���Ie1�Ekc	.�ȣF���Z���ٓ�O7�X�-RR�����	�3M��{NI��!�m���7/p_Х��� G��\�i�0D�#�m�ټp�0�_}��a�;�i����e4C�T��7����J��e�qU���ۅ �l((%p^x�KΞ���,"1�a��Qu�Z�XbNm9���H�:]:j2�D>DO&]�@�-�莒I�J8�,���eL/�~�ͣ��1�ɻ@�o��r�O,���>�N_E��a�?��?]% S�0** ˪��ni��䅠��ԏ�79�c��L��Ϟ;�2s
�$�۬=V$��0ZCM����.�J\�8�%8�R{,��8+F�w��(?�7KNG�k3�qx��Cu�Qv��ڔ^M���0ʸ�U�H�J�u�� Q�U�A���N��ѓL%���f�k����b�K2Ū�Պ�:��o�	���mS��Lv�՞Q*�s��hjVkf��T�M��l��Y�f.�t��A��z��T��S�Б��`�����e#��S�w��R��O��%l��T��E���3[�pXO��0�P�X���9�(Ġ}X t9���*ǲ�\ [��9�8�T�V��ɒ�q��]�,��|$]��|j+�.j��l.n��s���֖~�R����"�"~����Qsm����
�Ӏ�(*DPx&+�����"�\���L&�s'T�@�ڕqje�����G�F��f}+2�56����n�I��Os��tC��4:���R�=7���B�F�{�$;���X�.]���-\�R�+>(�,���C��r�Q�D&����`��& ��� ��Wd½|��;>Y�ؿ���`��c^��חY	Er0t��G%K2��vt*��0F��9vɽ`W�Fy_��*⻼��� ٦����(f �싐��q2���)�7SA}q���'0^z��>��a��eaݾ����� _��.��;Lh�V?� m��o8(�Ia݇���v�"}R�B�57�S��e=�媆�ƴ$�,���	9�C>݁Q&�G�F�IzO��6�W`6
���:5iY��P]��ĭ.QD���y�f��_�>7g��2U�ɠ�ea�iN�!<���^��aC�Z<+\���[��U�B3���l��({S����DJ ��t�qV�	d�U&�k8<%��_.W�������O��r�n�KZ��T<r�c�����+]�"l��͖I�]w�o��vy�ީ(����׋P��Ż+�����1�7#G&_T2��
d�hJᢝ\�r�-
/����	5^��V󄤃q����=F��Wa#��!h���|��,r�=���]��ug���&3�!<�<�_nǷ����pTx�rfj-64�}�������Pʷ��obU�U_!'��Q���/D���ҳ��A�C�d�鬬�j�~e�����L�հWg�#�Jn���4��3�NJ����g�@r?9����$�,�Z^�rQ���QaY��宰�G�}���Q ?A%�p��D�LN�=���JC
E�ѕa3Hd��(`+��`{fA��)В�I�sIs��Q%�F��[-[ ����!�Q��$(E���v�n�"���Iq��ĮcM]�����;m�T�\q�X�L��F���P����b��_�ڃ@��S�k�+�x�=�ݕ�X��)9Jr�䦩y��-obp�۬�&t��l�kH���>���?O���~������7��S�����"�.OW+r#��Z��8�z�Zy����
�k�Sq,|N�C���p|ZD���Q����YJ�^n�i��	[�Ty�9�C�Y(fRsx3���d��������'ʎ���X�T�o�5����h�ص�(��оM*��!�WÜ���g[�A�cX���X^����Z(�6J�����S��M�*�{Y'T0��M���%�ו#
�s��6�cf�}��H�L�����������lS�\���I��Xg�X�� ����Dk�*�)"1��^��D�-�z��.k��@;P��:B�����cGX�h3ާ{ X�� ���i�� ��#�JĞ��E9�VJ�m���DN�^3�o!+�aD�48�C���%9����K����8�u���8*��T�>��I�K���Ό+C����#�o����>o�2�X{����}�Fu���W�!�?�x*P		��?W�6�\�xШr+�6��;;ڒ{cG�^�=L�{�C��G�7�8���Rw�(Cy{A�pO�>J��Co�ˎ_�9�- I�8Y��z��AU@�o���o���F�L$�R��	��wI�[A
�=�����5��h��C
�'��T�W��$/91˭�e]}�?h�e�oLr�rBt�U�H�0˘U��ّ�&ѿC,�VߝX1���]h��W�� �k�`���ف���|ܖ%s\��R,��iP�ld���=M$��"����^r������%T꘣Il��޻�pݺeG�FrN[���܇}����I�>�`F��@� L���y��	�ij�O+���Cv��\�`��[����#k,��K�����`���-��|�ڂ�1�#2Ⲽ�^��)d��)����"���ƬZ�xt{�֔y�B�*��V҇�����H�dmU� �1�%B�wI�~��Wΐ�Nn�A���/侏�'�v���6�j��W`�A C[�z��1�]��b��a+�7r�pϭfeC���ڎ�6_�XQ������_i��4��~'5�P�����A9�s7v��@��4���X�����|���-x���z�ԋʊ���Ħ�^�v�	�:n����W��*� ~����Кu� ����\�_Y�1���:�-��$���D�'}���u{�w��y�蕟à(�v�Dw觥�dn�`	�\�IڸG��p�������,T��u4��\t���:N�����pkG�H��Yl"M�H�$޻k2�e��J����ܐn��'���������8�\�M��w��������ŗX?T7Ag�]�%�@`���'���N���9���v"�m���U��J�/0���CH4�a��Vy������� ��I�}�ݭ��Š���JS�dԖfgm�r �>Q*�	��[�>^�8Iv�s�;۠�aA�_eͪ4�X�E&��Uv��W��{��yak�!G�!����Gݾ��v���O�
�c��"��_��@:Q����ù�Λ�x�K�����Yk(��;p��D^ɖ�m�r�gv��:�>^M��#���nrnd�]��ڬ�����Q��O�qw���N��R���?UP���>+��o�ڋ����OM��?�r�|���Dhy�L��1���A�^�.%|0�I�X�%B�&�eOǵ9��U�K���^QM�7�W��A��ܠn���"��CQ�}$�)q��o|� Dc���]���Ħ	��藵�o;�.e����GY�|v�J�� ���A?��	_�S���;A�h9�KL���aBl��_�W�]9-���ϊ=Ї�Nv��-�B�E�o˰�y��'�kԜ���u+��._�G��
�)�F��)K�W��'v[ƙ�6���z+5�q;�������
@�c�K�0�-5�v0h��'��O3JN_�N��/C.�D�St�}�<�ú8�SU��/������|�`�Л����l���k	�*���w�7���ؒ��95,�>:�W�f���-�;z$<i�0� �B��R����$�R
�!���ye��@=I�U�� �En��k�oN؉�T�K�_:�ӗ~��*@��b��7���0$i�	$���#6\4����/��"[++k�i� �Co����_�{Q3����m2�������bG-3�)�ԫ|�yoEL<?�7EjݺmAE~�� �5��v(V[\,m#�z�~e=L} ��ڎ�G��	�)k4Q�HK�P�t4��TK�[�>�t:��shS�UD#��:_�3����C���83P���J[C`;����τ���.�S<��H^*�N$r��z��-��ѵ�Y.�n^AaEΟ/T��M�_�h��4{��R��==
e>Or�$��b8,a0K��j4��X]�L���F�(���*Z�#`s�ɬ�6K)(��i����Ɏ���+R[e�ϊ��݆G�zJ��=t�-8�l��c��:2LR��tp�Y��p�mc�3ܖް0j���m!���P1�'Vs�Bl%O��0��!����A1ۚ�Z��ip5Wa�BG�����w����
����-�!��Ũ���Ɔ����L�Y�H�Թ�S�'�~eE[���C/$��T��<U\~��X�?��%��L6�l�e[�Z�B)8��ecuFIoq��\�Z�7���d,�9�`��l�Ʀ��Ddui�Ե�bX*b��?<y(��b-
U��Yr	���P�����/�5O"��7����_��3�0�G*����b�8{����CX(�B���dBK"��Q-y�@X�s��F]U�%b`���G}��V�"�'VP&��S�^�*HWNyXa�9����xܞ(���˩I��/∛X�/7�S@�b'J��M��I뙫7�Z�r+�0d����0����0�R�<����OAe���� ����w�@�t�.�����|�n�[��95�"S�np)�abs�Z��=GJ�QƜ�i�:�֫���\�/���1�r�^�P�Lb?2�*�h7ZM-�u-�|����!L�B�`�"����Z�z�H�$�R"*�7����16���(�P����.��"����hԀ�5F$��.��2���C��냶V��w����p~f�i�9S�8�U���܂%�
äG^�?���LK�uN���NM���V�NKa������n���u�i3M=�����@����N�����Dy�nR�t���nj�c�����Uc�9��dHa�F���w�:�}��4聯��`�]<�����9l�R�D�O4Ws� f}��ԙ�)���L�`��2�@[琐�O(p��E��)��5�U 01&�0p�lT��!I�@��8�-g@��!N���-�T���t�1!��!�e {�'�ȗ�ӫ�dr
񤞲��0'��d}�n�b�t	��ѹ�a��R�S{�l����<����~�ɓ���B�l�tؖ����H���a�*7�̵NNg;Я��cc[(�#!�Mu¥���#�lؓs�]I���ttH=��^O�]-�y"��rW`���7Kn1���V�Z�3����V�
]�����*����N��%�r�(M�c�RFM���R��iG��_Db!sͪe���ѝ�<RG���kV,V�3A�w����(>�*w��u��kq3����!#v)"������uo�AV\�9Q�c���3q��\�5/ë��p��*J���b,D:9W9�8�ï~k���Zn�|�|y��M��5��g�5���x� ��|˯�Tf[��˃�����;�������`��ݑ�",ܶy�Fh��?ڲ�	0Z��o鈵[�Mo�B2���Kt����S=�:���8�/�_�{��b���A����u�|�����?�B�먰��@2��]�N�lk�MQ�@�U��h�q�L!7��k	g��W(��l��~ky����/O��u��@�η�[�U?a��oT��(�O%�z�5|Yi@�vXؤ�bx���P�š��<?it�5�;I��8Z���������XKZevܑӁ�ƩB��VSBN� ��'�C5E�a"�Y�ُA�5H�����I������f��)�<E}a��#'_�k�^.勍C�d4��}�ڹ�,sV6����t�Γe#���{����� ?@��JjJG�U���>�9�;kE�Q+�v� Q��Ŗ�)1F�]{��m#�ȶIX��S<⧖ UQ[2 �n�v�l�U��:�M$]D�3W����?���.�Q;������+tp�zA�Q���]0}�"�o�d߁-_A|��s����Z� k�3ëZ�h9�t���R��c�w��8�yj�6��U�:%����qvأ��c��{ ���f&��
������sx3�#��4����;�$^:����4ADW[��ǖ0�`�;C��[�`z��A�x���61oxQ��%ꍡ|q�7`��R��u �ѭo��8�����ƙ���mV���8�H=�ͭt�)��������6\X��/��t<ԍ���o��U@Yqݶ|Z�  +�h2x���1�4�ۋ�s�2��q�!���� :)��_H�4�K}v���N�3���8u�����[�d�kD����&S�#�Ai�4� <�!EN��V@��s1<:7�4?`8�Ȝ�ЁL�Ób�t�� �$n)�A�&�9��ՠ5(��ׄ�D�c� yZ%Ȃ�Gi��FZ��j�������a�7���pD�Y�E [��k�����r	�z$3t�ߡ�t?n�*Z�V��5� *��hZ�]i����W�CBf V5W���������}3/��}8���P��z4�R�/�G����[���6�ŷ�ݎ+ӈ8Kg��S����.ⲱͭI�l7a�Q�k�,�gZ��=�I�F����:��]���@�s~C� \�∗��,�ى�ꢯ��\sW �������ե�OXL�d2x$Җ��rSV
��Of��8��uC�V)��#ii�w W�nt7u���=c��vz���_�pX��yye0?b/���d�p_�@�������q�m!���y`��k�7�63�)�����%�]��>O	�ķ�ݞ��3��$�uŇlI�}P�7���-@g�<-?'v�����٩�1�J���s'>�7k�Ȗ�=�'�2ˡ;�\�N�3���e�y�ñ;����~��;��TM�� \�̣��U\����Rm��l\:W�-�(� \���;=�/p��o���Iu���i��H��랠2hܺ.5UK}����٬��o2�%�t�#|�d\�bj�{�.�!�9(��on�q�}��O���*�lq,>�!�w�P,OE<��=�V_��c.�#�Y�}�{K�	Z�7&����|k��V�-�iN�]��Wq������G#��j�*W�M/��m��5u7=<�b{�|ݎ�5�E`�A���M��d_�3����^�
�ah}	�vFDL�F��0�����v���xf!͊��RAP��j�'ݵRY)�
ڐ���s���u��iuq/�`a[|s��`q�C��:D����#�bFN|��y?���?u�o���%���ً �A�V�Np��cF��x9J�΋�I�j��d�l��,ȇ�pg'C��F�m]/X� KM���&�M�֦��*MvFN��&��i@p�	�4��!�a�Gݾ�8ێ2�|o7x�PmR�#����p�K���~n�	yt��hlj#�2(�����'��t��<8,e���\��0�Z�;����FCU�[ ���%���r".d��>�w�����Pf�XSW �%�������Df�t�1Si�l��&y'���gϤJA�L����F��m2(#�ZN�`�Y�xw"!�Y��
��S��L]���q���q���E#[�T��s�	��3�*�p�(�8b{�Q�NSR#��Js�H�Q&�p����s�Q���=��5]���4���&����e�� �Fk孷ō���R�)�B�rc2��d�n����J�kԴ�Nhw�
2r�7�Cl�Ĳ���TC�� �3
��� ����jQ2�rq�
�t��r&`��C����h�I7n6�i�Ւ1��6`~I0�<9��y�N��(n�gY~��	7��5�~/8�������͍��"��/�e�ʱ�ul�����'`�s����'ED��wN�V�`�j��s��~�<�0�"#�+��i"-%`����B�����b,u �$5Ul˙��ҧI�.����X�V9�=W�hR�ݻ:;��2ȹ�r�J�����t9��/������k�~b6K�FƗ�/�&I��\��Nj��%��a�%gc8��� v˓0,q����k�)���X���$���(���<>�x����zn`�`��"X��gݱ�8&-��׸
=��1��F*B}���S�2�:�
,�ޞ0>�=M�1�8�����d��vs��0����ery��Q�e<�8k����۩�b���t����̌nC��yսA"72�6[&�\���?���B3���Dż��!F�O"1�N,�|�����I�8�Dv������η4����-P(0^���Щ>�҅�Ov�v�}��ˑ}�=�
�q`-ؼ)������;{e�J�˸m|e</b��2 ��TԤٔ�o�$p?�߄ަ���9g��L��*��VS��e��4��J@α�h�!���2S�V(�������g)��H:F��Cc2s���.�P�i��1c��V���Fǖ� v��Q&?�����hׁ�m�g;�)e�>�$c��5v���ho�
o��2���jUׅ�`�釽�ݥ]�[�����eq��v��$E�d̓��n�0�j���Y%�b�UBF���<� ��M�jRt�_�x� `|��z�}W�+��f}#�>��-+�ȧ�W$2��w���O�12��zB*U��u�H�nz�/�~=�y7����̿�w�j�#\�hr��$.FQ�rٴj��j�'|������/4�g���K9��:ة���1ڝx�����]m��M��ヸר֑lF���=�{iyINS�9�����.w�LU���O Fc��t��CIҌї��@uui�\��? ���\03F�����S���qu|]�;9}X�q������7�BÕ"�o�b���e�������\��`�����<_V�G͹B�xnJL!���[��.e��9!
W�/_�����)�|������ˍ�)��"�<#~p��+�6�ˊ�ѵ�ű?��A��JD�V$^�T*�,[RH�ȱ)��w&-h|��'1 N����;P��i����֘rC�O�2��ɈuF�w!�@`���˗�@���6�7��j���7��;�e�TW��h���f棚����m7{-~��	(�\��:{=P! #�h��v���-\��c+`�c��v�H�+Ɠl~��0
�����_�:�W}�ɽYF5�UNPV<�6=��w��u��qn��Ē=�W?�U�z�"�.T�g�ڱ�&W�|��L���H���K��p��ޮ�Tt�����b�T��YȤ�@����Wc��(��ED����3���6���Hj���}�9��A'�#�XB	n����N��<(�S�:1�/��ي����5-4��9Ԉ�R;�m�N���}#?m�"bUg����_ua9
�7\H]q�^At�����pQ�����I9~��u�0.��$>�`\Ln��9H�LA���hr˂�k�A�g?X��lktL�u�sU[� H0O���pR_��BȚ"� 7�u�+��&�PZ�D�JcZ+SIS�O׍�I_h�