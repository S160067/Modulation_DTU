��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����>�S��fI#�l7x%���$or�#�6�y���N�i� �D��f(�:eǊ�` ��S���^�mBƱYjA���v�0��kh������#�v�(#W��ux��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ�A�O�c9b��2���j�:��HA��?�\/��q�k��#W_�0����J杦�&���£mj��̟鬶�Pf�s5��q�Җh.�k�/��HJGS!]$�y�}�t+��`O�u�_|U�� ��4Uy�J��@�h������ �|�.��oc4��ܘ���xB�s^'��Yt4�c������~?1�r�ȶ9 �����o2�g�Ck���%�����'1���CE�p�X#R��(�Y�6D�p��\v��p{��a�@��t_]��j'CfjE{
�Q�"���ڳ��?Z؏Ζxv ��n�wg�N?OWǖd�0�͛�H%�}�B{�J��yn(��ZW�����n��[M��Y�@�p:U0_#�e<����O)<�:8'4�}� �vOW�%Œ�C������*��ۭA�f��>1�;o�����#1d�3�J8�*w��K�d.�N����Z�k��(Z�#ϝ+ yO
�����r-��5���ʁ���SD��?�MA�����^�%����L����Ö�=#���Vxgו4H��J�.UR��3z~ZY�:�c/�Mw4W���X/�"s9�nx��W���7�0V$j&��[��ИH'%c��w&��v8�gm��=��TB���[���['`���^�9��TN�m���,�X����ո��G(�j����3"�>�.���:����7Qޭ@H�F�=�=�K�#�Vm���^�	�o�LCR��e���b���٥�:�#��I�SXL�,d�9KIM	�P����Ɩ����}�<)f7[�{�l������ȓ?v�ռ�_7�"���pSJ�:��6�8p�v�_��I-E��(�9-M���0_`����phʊ[2����?B�?�������3h�O�I�$�H���s.��L�H��D6/nR��P����|�H��������k�%=j����?b/�.��[r�|���	TNy��F�Y���Os��p�(*�Abe�Mu��qSV��m���F%Xl;f#�"�a�Yp! q�����r�_��G1�qf��qз�h�a�?�P�=O���*�v2 z#FH��p�-6�t�y^���D��_��V�O��8ז���CQ�p�ty�����U
���w�D˴&pR����I\�����N�dzU��J��f��	/i��5�'�Pؑ�Cf*���QM��]Y�B_��~QD��^������fё�r�Ov�H,�.���;�^EV��R�	���H��!ƭ�6��-?RvV�����0��&Q�F̋�<����ː���8�;�#�Xa�� ���~���A'����E^�$t��>����[
�����lQD:lT���P��EMt�E��wn=�6�'�S�D���r�,=����|�B���q夓�+(����3^w�?/L"�E����q��t�$�~���?K�No�K;�3�17�3sv������NJ-�y��h�54/:��AU�{�p@�s5z����x̶�{��vK��r,H��qA\5�'�z��N�����W�f���7ex��E�Q��y�K�pkQ�2GRd�L+m�����4!��rd(��z06����p�h�b�dF����  ��Ll���O��E'�!p�Wf��8���o�/;D\��^
F|>` ���BCe� Ry��r�w��0�v�t2�z�ڊ�7z�|���9��
0��O>K9G)]*�8qv���H�ed'�bJ"������ﾷ�^�*˲OԾV��M׀B��H���]֥�ԇC)�U�'S�F�@�$_h�?m/?��Z0���^?L��u�N.��k�<�k���'��,��Έ�'�Q�K���q���8J�= 頦
�%2L����w��p����Z$�,gNkX���C�����[%�[:D$��ͽ�g�Ο0���/,zxm�ޞ�Ce�,��Q\N0�YI��{){��D��T�q��|*�B�tXE��p)�%C���ET����kx=��-H~2�~n��t��˽�8������[u�� ����X��,@�V[|ztO�	H����`ן��+�y}���V*6��$���n�d�k���%3:2$O{��������g���b4g|�f��
i���*��<����Q_�s���)l���O?J'ؑ�m��0de�d_'�k�(���Ws��EϏ$�3E)�u9����~:d�R��?G�Y(1��k�H�.���X�cJ�@2+d�N8�S7l:�^���j��.��	��C�:��f��`� �q�ٰ�� �hVЏsB�,��D�'����cR Ɉ�fAg�{A��P�fC�x��<R���"h��A^�!Y��Mzv"s���ƨ��29ބt���R�D��t�E�F�ᇚ	��i����C<��G[Ü�l��v��OIy��Z0U[�a������7�F/P�izu�{7l�Y��*xS����z�+Q=7;��!��Iī$�y��뜰�Y"e3�	���#�>9~��\K��id�#]��=�]�M���s����;ui�U:_i���qF���5��ʥ��"T_G���)���j*C���IRN#'���)�_�;�~"�3��a֓\$]�I=��`[�v���8D�l�f]}x�/�lv�+X�o7eކ�YMaIX��f����
)a����e`Ƙ(�Fu��ׄJ"X��t�.�-�Ƴ@��!���kZu~���hD��>v��J}��`�ţP����Q��܈��xb�>S�����V�30�a��!�`U-�-�4�R@��;�N��]�Ɯ@�K:�fTC$���%)+�v~7&w��§̀)�D�i���m��꤇��}�o`�n,'��%t��~i���񆼭;��o?���P�@����x��EF���m2��f<*zf�����d�kJ&�p����"8zWxF�w����c'0.`��#��i�-�T��ǓM
j�鷍�D�q%��I/\���VQՇQj��6�_tf�O	l�U#l��?�{P}(+|�7A<�	��.OՀ��Qs辏W��K��F�5����횶�`�V��zY��D1��<���2x��/F��І�@�,H���؁��$^����Y80�]�@d�Z�� �'����G6Qɼ�1 �Pt�^a��bM���V`:5�H�B�\_/���G�jS>�p��:���w-����
r�^&-���m���\��ۆv��+3�8#�qh����se0)�M �)S�Tw��}���=��|j����Ev��[��]7N��]e�{6����� ;l)���Zn�n�����3a$�ɱ*�� oz��e�̙�~�Ä[1�(���ϛ�j	�MXE�((9۠R����IF{���\�	��l�8.�W�� I�;َErO5"�.��d�V�X^y~T�<���]�K=dy<���V��$�s5�hI淅�.���>��s���zB��0����X�+Y2_�5��K��x�i�v �!	��sg �����
	��D��|(��"83�� ��^gЇ�p�Ub%֎1�5��&�k
0@I&G�e�G���~�?͔��+�_X�\��t�=1��Z�UR�Y^c���
���j���i�W�Z�7�z�(������ ��<����@[T�M` ��Z����<�)�5/�rm���1���+K���B�z]����_����Q�� ���N�v��E9w5tV��p<@ +vU�$��>E��P(��|u�� ��h��������18��	���]��B"��U�f5�|boa������f%9߼����$�/����M�DGT��T�w!43Y��Xe��Z-	�װ��>~D���ƈg�c�����8HZ��%�I��6�A�G�ګ* �� �JD�y.�y��q���'D%�8���͝BQW����u��d���կҬ��i�b,3�(W��#��{�-]�����m���u�)?�ЅyR�1�Bջd8{g�O7T����N*emL�&h� j ٵ���Z����P�_X1��Jc�=!��x��=贤�T
�`n����p9s&��2$ E.?`�Hm�!�_Ձ�-y��0�7h+�9�)��A�uT H[���p�6G�<���n���[ﮇ�ukr�r�]�X&�QBPu�:��(H		������z���bAΣ�G�����m��]����os�IO>'��5���Bu<��4�c�X?s�x�����*���i�z�9�(A�ؤ])W
�<h��m���x�V|7�C�<O����ii*J���<ǚBcԌ3͘4�D���eiHښ����&B���D<���!"�Cz
7��v.�����O�`�o�`L��E7�C���JD3B,���g^8�u,��4���<���`TO�H�
A�?�I8( Y��d܄d��+䉧s<�|����8�Pz�ܴb q��Q'�=@5���Zx��$���f�@sOԄ��v�g�@����k��H�rV1\;�Š�̓a���Xpx���s��7�����H�BG���I��t^��#D6k��:��#9�U��]��p����
�lY�7�&̰��[T`�֥G���CY؈���s�Źe��ٙ�U����w�6�h�N�^���|�&Zo�h�����<W7�L����4	HƯ-������\�% ��u�iLl�^2u��\����[��5��D�w\-AC4P �0bg���k����^}tݣ���u��V����c�覣��1��=��_t�&`�oѦ�'U��E��t_��d)�N�aP `ωk��Z)Z�rS��TBY!RL�y�w��F�\�,z!s��o�"���-� �G� L�X�i1����L���b%M�%HY�a�ph,��1<�J�c�2��Ύ-"7P>d�b����t�9�T8 �t{G�P����r��U'��{O����e�1��7�_3���M�Y��eEJ�G����1�Z����	��S��Yͫ�
�tȿ)��%���
��*�>5>�֙�(W�Y"�7�$)-���n�ߗ'���b+�>��0MF¬*3U?Qr�;;]�;v�ޠ�Y�F2�ы���wI��[��+�]`&:�;'5I>��|���t������>�T�t1�A���D�F����M{ً.	J�!=Em�?S_��W��c&gu,�.�D&y�(�]t�d_���)C���%���C�E3� []���,�(��miqKK.���w�s ATCK�AQ��򐭊�;�.�˧�.��*���/$��L{���ʚE�}Ep�&F��O�...b|u�R7;τ�=@A�n_��Se�[x�y�n��.fY*(?���%#�0�]�OL=Q���U��w9�����2
�N?N���ȴ�@�>[uz�!�Qcc�c$��z��t�_c#.��̳� ��8��]�`�����-��'a-�A���vQ��@ff�/��"�0�-�O^�dѕjSꏎ���'��LCҠ���<H�<غ�>��Z����~��ze�:v_��߸KYa2�K^eG�ʳ��@о�,�+�ͪ��DYE�����(�`Ԕ��O$_�p/	a�.~���A`�fX7��}��m_����^LL$��o04��Ol�&WfI��ph�N�cxl��w>Z��kW����е��8����^}�@����	g�T��Yfu&I��}��2%���j:S�4Xr��>v�zR��νPj��k'��.>�ۏ6M5F�j �`L�Ԇr�B�u*��$���N���6QzVW��9��������L�mni�<�zMя��6��FJ@ �o��B���Ad���[�;��K%�i���J�����aٗzO�0iO,�ӽ��ĝ�i�

9�r�~��=���r��wE]���k4�mM��û��hx�D��UǍ3P/�T��R^_k'�Sb������,�Y�*(�y,i"�p:�_6��ҭ�dl��op��z2&b~�*_46�M(�7K�7J^��ȱ�(3��J�+<�g��4��Yg�l�l�nt�H�+_�`��"�v`�(h�ףS���ݿ�V�9O;�(P�_��Y��5�>�ޘ�|WDuUc�O�^�Q������>�
z�:��TE�Pi¬GK�g!�^��}�����q)�+�_��3 V8�N����TxE[����5+
k�j-������=ל[�����*�GjW���x���
uR�L;��SGe��;
�ʱ�3������&OҐ��vw�\q�m�Zq�g�8q,�)�o���K��]�3 �BN��0���Pzy�P�\�=����a"�PẳK���jP��@ �*A���ñ����9���wY_�M�=ў�0�^�֚c�F;��A�Ǚ-W�ET����	b��]��m�U�*���`�h�!P�M��)�\ɹ�q=�,[~�D���7,���cg�>���HN��=bhGf�\%����Q����ﱎ�W��Fa��}��p��~v�*���=Aa��d��iM���6F7�-��e�A���m����A�	�8�n|��F�JQ�O�+$f��o)Xz�*�9��f[t�]@i�|8'�0�y����j[�9����:L��S��IZkc`H�O�>y��y��( �Cg��Zխ��A�����T���U +����X�f����Z}ф;�i�<��Mƴ]����Ч~m��� =N��	VB�ht�����-�ڏ�{:Km�7�K1�c�YX���vz�U��W�@��]�І�f=��Ԡ�L�`:�3��oUN]&�a*0ѡ0�w�;�g�n����/)^A�� �\�r%IjTT`Df�d���=�F]���M�3�������T����r;�ԕ\,���ɸ�I��f�Z�A��C̵���p؇�u�B�������3B?�rx�Z���T�a��7���$��}����aN{޺&����_���}�����C��zd�P�ȍ.�E��B�`�>^�}��-2���0~�oH�}���Ī,�yl���;g����V�)?�o�|ባ<
?�R�[�}������ޤ��z?6O|t�9�{���W�ꭄ\ ��}I�.�C��	fcr��,��2%��tSJ�k�:9ے�W�a&R�o!�ŗ���m�ئ��΍J���0B�B����\�@ :�p�p8U�Eg�4��u	�+u�OmdQ�R��X�a!`c+���C9�,�� �ں�-1��R�M�
����G�T`�?�Sl���/�]tn\��D��?�ړ�G�';p�i����F{S�)��2��-Hd���ˊvqu臸B��ӧl{�$DNu��&�Fz�m��K9KIRF��y���</h����K�d���,�tiN�z�~8���՘ׯ\d;=����1RS3r���l{�A�#XZ�Ӥ�N�Y�	x�H�1X���ss����eC��ĝ#�j!��da�u�F7�p� C����[y��u�|�͕�8nfI�Տ5�v�\��y[8&��j����+*�v�_Xw^��q@�S�S	���\���L�vO0������%/���ܭ��e&�^ �^&�y,M�0���RE�Z��y4H��/3H��4����4{�pz��.��.vgL̮�2��pb�����g��]���W�]��c���ԉgjു�[Դ;���7��lS`!�(ƈ'�z�\QY�1�5��Q7*��-������O��_�-G�/C<�pERLhE��f�Օ�� zw��SU&tb���Գ��\?�E�čӏf�������I���+�w������y|�J��bj@zUP}�3��v���<�!(��?B㒥���5�>�z|c��(a�_��K;U3��}LG�T��&^���(ӆ�s>^�4����8^AYG���l��qNJ�x�	I�'!���a���Y��1[y?�l�'��]�.�dgћ�zZXԑn�LT���s&U�H�*"��}�Jh�?�U�}�a�������V)%�hL-#��������X��q�}�Ͻ
���g��)�ǹ��կu	�a%
��I�Z�ݟ0�ƄBln�8���,'�C%�w!�9���K��J�h�����A���]����t�j�s����}l@���P��VW�[����T���H5�>�d��F�G� |��ɱkƤI}VM?�2��((VS ���S�/����~^?-St�n�CD}#�|X.�ON�Ul�o��V{	F
:�\<�����>d���m��뾸��+��8:Ǚ��A�W��.�HF]��a	�dE��[�Gޑ�W�ZV+�/��.U΢����t��$�:�x���v����Nb�6�y� ��a��&��8v�a���s���'�&�q�̳-|h��Í�%��Yp����bӕѶ[Dlf�:�`��+)���ܲ���$�Q̙��K��c-�Z<5�.+���zb��ű=S���#y�8\�m��Y�DaK������8X��Cڧ��_M�8	t�u��.���4�U?_�-����q+��ƕ�iϣ�B}�G䤝�.����+���F-@�	P�B����>;+��,S�]��/��2�m[c_��s�K҅+9Si��o|��KU9����[;��9�e���o��x����;Z0T����{O\�Y7y�3�(4�sK��y�2϶��yxJu^I4�<%"�ң�M�F��(��fC��<�V�% שd�{�Oҹ�~�1�����?%�ET�j
��_�ӈ�/�t������P/��GF�ٗjE7|�k0�?�$˳"}u���+�h�f�R�E�E�W2kzۆ
sW+����x��)�K�X8>�'�J���g�����\T!&ϐ�I[�;�/��ٞG�;�^����Y�Ý{_��|2!S�Y�1Q-� �m���"8���Y�C��
཰$�6�C�Il�Ja;�����xҨ;�G--�����NIáW��)�����bu�������G/eV�kD@z����np�S�H<���M�/��,T���^�>M�;$��^59�
���6�nӂe���e
���h��"3 ��ܴS5�6��=�,5��[)�/_d=���7��
o��W;��G>-٤#��qn7m@ l�-!�=���#�5��4n]%�oQo'X�"��źF9����^4�hu�@��S��z�vPoC�)
n����Nq�,��t�Y���W�,�۔�:��0�1*"q	Ms����iAunTN����g��*#����Э���nv��-/�0�:��mm'Q�`��X(1���� >a��.�EY�kW�����;���A/3L߮��-�S;���Ki]>���-�&4��T�/�@/�ej�Bbc�< (;���	�����]��.z����/��P���!J���+�τ�3K:.g�T��!�l��M�T�WÖ���Q���S^)�n�~�����݁���~��uT���3B!:]�ԕ^�2M
x0�%mϥB�V�|��0���\>^Lw#L�6�i2Z���F\NU"�@��u�F�q�z`�3v�l9��ʇDA>�Z��Ճ@uDCi��`�}����ݭ�c��r	�S����w�(���˗�Rs�f�FL"�����on�����	A�f�h�*D����(pGH�H�l8�hz(	��H�n�$�DJbC~ B{/�7���Ct'ܳr`<[�ȷ"Ù�G����8���&��K��n�~��_JqM�8����T���=I^].��U���_fY���/����5T�e�Gf��]S�S%���5(�����,�M�{�V1"#m�%E�!�|?]�%,��,_>�Of�*��'w�9l"s^�,�l�L�1O���z���$U�e"edP�#bE��џ���@�G�w̊��R��`&��1eG�q�b6q
�C�Y���?���ѶT��F6�65"�߲�����k9�[������W|}o�ւ�rE��d��;�7y��7����3����Wln�������������4��u��Y�ǚˬ�PD�ݽ�\�V��4��O�����ե�gͼ��>3��!�#A��q�Wk$��B_ܵ��^�=q��[:�8\k���a�e��ɮ*V��9 ˳������r���`���)F��L����v5H���G��(X�<�i�C�{1�E���9Z�G����h4E	>˝U{�5��c��;j�VȔ�D�,�P�W��o8;ϫ5������T+"����/�by~,9�k��ԄޙRM_�������¤���^��$�*1R"��5��qT	u�/�p���&�n�G�l���Y,�ܞw��������O?��Y*��O�yL:-�= 2�S���/���r���ίNq_�/�ʑ��ÔfK��K���,�����p8�V��
�����SU�60Dք�9�AyÁzY���m���,������vԆ<>�&�rJVM�YlT���ܔ#Q�ߟD\���>;HG
I�
mH�7:�l>^����Q�"V)�ۇҒU3��?��(u���ᗳ��MG�:�8��L<��+5�݆H�X�㢢j��S�^���>nZVۼU�,x`���ЪB���]�ܓvϔ[�Q3�X�/ú	#��~��%۟��"��B
�O�k9ߑ���0������fޅ53{��{Px�qW6��
���y��ҟi �b���JR*@jX��$�y� o�>��, 1��7��y��.����L���"��\��dR�d	��H�����,T�"�%t]�<pE��x���װ:��b��Ze�Q���B0��5�e
��s�RC-�;�`�/V
+������`9}t����GOi�������k�Z�����q�� w�c?�d��Ҝzb��/�)NV�K�4?��AU1�� �J�V�;�fے0F�ĴW�dYc����A?���W�a�/*�F����U3��
s�T�w-�誮X!Z#�
��G�� ⏴��m�C�K�!I�e���wkf')P����N�'~�3��o��.5aB�;KL�fO���u��)�-���Y/��ˋ�N�X��A74�"T�+�9