��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����0� ����遼�6������"���#�{A���'j�Qj} �}xT	g��F����a��f��洜K%g==�Z���L1������bG����XB�k6T��w+F��3r1#�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�O)E��ik�9q��~�Lb��,�J{
�B��Y��7�I�'t��qc��^��	TJ���#�3�"��d&�&�{d=[�x��krWчe�>@�h�3M��X�������f���<-�TLTe񜴦O<b�d��#҉�6}j�h�^�6�U�͗_�u�)�(T��4���H��qu}GgM=ū}��}]i6�cZ|D'&�+� pe�H1p*+��(+�c��ś��è��\L�o5���<d�v�'E�B㉵���txY��y}���ȫ~���Zi�V`�4��}��J��V(&��y�'�u%�Pp'�� _�x�ƙ%Q��
r��TK��!��P^d[M��لa�e�vj,]ia�)SIn&_� �иb�]�+��W���o�O'���w���i"�In�"ąR�'�?�]T�6�ș��m�!����j�0Nw�������w+g��z�||��6pEn�qƵ���ǁ��
�Q�t��?�2䕰j7dAL	G�)�f���5^��x����:I6B�+?ħ�v&�U׊�ڎ*j�|��HO�E�@Hf[%��[>�=c�+d�%=����{�4u-��J��R��ᅋ��
!,����^���{~���VՆ����0�?u�k�V�T��8)ŏta�DV���[��lF�=
g����w�e��3<�|��6�{��y;��EPN�'�^�$��kỺ�M˯)�P��U~�Ww�j[�c�@���7�L�����#����P�t{|x�ا���X�DfW�~��}�����+�|G���h�֙�}'O���-��ƻ3����:.,LI�n�!=�N!��&Sy�8��ɜ����"$�i��E}�ϛ��'Z57{�_�i��h��'��(�.S�(A�5(lg��>�����ΐ��B�|{ۏ�K�H��-Y��_.1Ϡ�����GP`�f�p�(��RD�2�������48֔��  {�.��-�M���1.���5���ϖ�.� S��3q�N�.�rP`��{�k(�*P���I�S�0F���J�8jZ�R.�1��l�sw2�(h)�'�-_F���� �h�R��Zc:�x�l��M������a��uW+|�j�����!����쭮NO^��
�P�W�E��W��T|��]��b�r��K�,���$��ݙt�0�����W����(c5G������H2p����{�T�P�u\\�b1�p�~1�^$�]G�6Xߝt{?K�LsQ���.��+�ϭ��1���-�ҁ���Qm��ޱ]���wG��-�F�`s`x�9·��̎�8�k#L�!�GxzT���v�2i�T����j�9p���c�5Lj*�As����ik!{{���-��#N�pD�o="��*��F��F��#S��#?x~��a*�mXz������>��(y�hʋ6���e'�]�t�	�2�ś�#�̳���axk��"{�#��2�&J���3R����^
1!��U�4�Q$�����+M��.�"*A�Lh15?6?kL�֠�|��]�:,�@t��h��ɆS�I��{?Zx ҄�N�<�d��;�D�ÿ�9�5��)�B�<�C�~���g�a*���L���n���z��g����v�ݒe4I=7���ª��sa�v�x�:&R�=B��!���5Z��S�hr���v��6cǄ&J?�y,�ά#��C�8�k�~B�:?�kjRv����[�K�� Ζ�~|�[��V	��� �%H����9L?U!��j�����(V�m�ɰmB�Aj;�uh�`#�6����=(�q~�@u]�){F$�3!j?[CF i�{+Ȁ�G5D�t��`
�*)�ͣG[�U��q�<4쳰�
4;�V�`_��,Cf�=�����Jm�e�UT���]ys*w�3}�S�(�ba�-K�q�>B#L��Hj�L��/�Ǆ�4�M��yʬ�_�Ҳ�:���Ƴ±,��>df����N.Fl��3��+*�=d� ����R�G����l�(�a���u�PW-�����9i��:�>��;�V6%�,SƔ)�jJEm�����`�q��6��/l�,4����2�0<$��0���<����3�kU<����]
c���b�\��2��M�ƚ3Gdޞ{���SE7F|RB$``X��w��	�O���n���u0�p���ww��4��= �␷�>�\���Z�97ep�hI����~�u����?�:��֒��R ܽ����v�q=�Q��9C��w�Ĵ��k�=ze�ῂ�pa	r�So��{(�$YSHs�0ו~�>�߾����Zn�I�61G�1��]{�gg*c+{ �|[\�a�+���ekT��J�Mک�s�P�ex�a3O��AWnي�1���W��#C��K͓��^.�3��)���TӞ����M����O�u��8hV+�o*������~S�G�8�+2��Zh�O��0�`�q�a��2����S@B��N�~���y�t�1��������䀤؄�L@p�lP\\3�#D�9n\����cmmp);f�����!�U�-+A�z��p㵒�ETt�8^M�P�L�{ ��>��,�9��,�߬����X�?5��z�y� ���ɍ�DY�Gs��?�U\˯�ERWD2�,������G{��o(��/�����5l��G^�P��5>ҩp���!0���Qs$~�>
�g/����J�e)7:��x�P�]}EA�+سd#	:���m�3�o ����pY�j�W�JÄdu��i'9Ī��5�%�?\���q�¹��ngA�$v�#D��ڏ�[D������ٺ\��pN�J j>TR�9�@��8��V�P�M��¯<>|����*��3  
���j� P�HGQ4k}��h_'�L1�uw[N��Ӵr-���OϟVM�I"�T��q���%�g��&�TA���M������F�+��.�CJ¾����}ML�9}��>W�6ǁv~�iɰ>�4�g�!�YX��1��G-r��lf���@�r��)�6L�g�|����FdP���O&�á�+;�q�L��.�|��S+�eW�\A����+���X�ܶ'�ՉW49h?�N�\�D.�,�*�a�t� 	����^H��^'J�Kť�\�pc:�V86�3B��t�;��i!R�X*�ǧw��s3]�t�ƧMH�ª�uK�
��t���\���!@#�F3�ۘf��C`x.7q��4L����7��2Y#���3D�*�Bף��ԕ ,�P;_�N�t�WRǎ3~.���m*T�T���w���l���s{�O��j�A�s��M�B�9;��A����8����'W$�fٹ�HpN�7�Dp�[��oH1W�Z�p��+e��۳�������/���}ԁLw�ڃ�ĩ]�i��G�3=�;^�P�6�Z�=Q`�d҈5�PD��P�r�&}�����ay�l����qK�t��a-�G���3���(M������Di�{�Z�E�[`f�Ј{�_f]�_���O�? �x��緖b��웍�����.�� C	RVA\G�L�GZD�?
���=&U5��"St�LC
E{��lo��*�*���0��3S�.#+� 	b�[�p�7$r�E�E��L�6|G/��5�e6x(�dӕSKu�v�!��ɓ�m��ˈ.&!�4���{��@�����`a�EC()���2���z_\YF(�@��׌}�j�Z�	�ywt��M_�Z�j7�6��_Q븐����o1���\):r�3x�$�q��U*G���~��SO�6ki�N�E�ʦ�l�m��f�O������i�J@��zX߉Vt�8��U����߻Dh����I����B��
f��E}7�s�EQA�@����9�������I����nD��l*y��"�]!FD���
YWb96~k��
���b�o/���x0+œ`ǰ��6����;w�Q�;ґ�h�9�_]���1n_�S!{��G=\�I�q�  �2O����� x��	���/�~�g�"5����޿�eP�` �z�\	ؾ)���}k3_b���3N.ܟY=�����y�J�(�^��!H��ů�F�7���GxLv�5f��XW$�Z�����@�e"�&e���"�C�z]��=���w��=4Q��db�6v�R���U,�~5L��׬i�.����/U��AB�XmO�iދ�$P����他���y�
\U\~����,�-I����N-q��E�Ri�tzHFsǌ�ۑ7�5��"'*5��ڊ~PX�@[�Dy{V�)/*��[z���.Z`r 
��P43]^.'o#u�N|�P���T�%�tCQ�3���W`�w�i�q~�>3��[9kU5�6��0	ހLL��I�$�@h%;��٩y���)L����r�8��~I7��u使�(�A�f��\F<����k>c�K�����T�)�m�Ýw!�o����!ꡝ�4��6���Dj6M���c�x&�15�"�* B`-��Kn6�B�ظl/�Vm�8Wp�ѱ)3��{�8�e�C|^�V&����w���7�}&��z4�Qr�+�C�x0�NC����&�>���\�V��Ԡ!��+�FH���_�ZU�6!�~���ʏ��K�vC�v]�fW%%%�N�P#|�p���\y���{GG[�#�0 �Z���ƴ�����ƚ�{
��]���J���w��e��M��a�m3RY��ѽV��RG�L�0��҅��c�J=� -�d3�;���C���9��A����i�zbyx��V�NLF��+PT7��а>�ŵ��\>��ɂ
�����ъ��[���4�g����~��J�����g(\{�dn�N��a�?����r����v���pe��4��K�}�"���}�@G�P��k��1B�u��=cT�u��&�ψ��@�NU�)�F*�t��r@ɯyc�Wk哞@	�ϣ�'A(-͂�D�ˏ.~
�-��(o!�%�(ۡL���><چ�������~Q�XϢ7v�Ş���^��)8��A��O|#����/��6�O탌�J�7Pe���z����z��ĩpdi}�"����S<R� ���!��!p��l FB\���Z��C��uJ_"IB�� E�����U2o�{= ��j��ݡ6��HnYI�J�Z�8#�%'��i���sf��N�	u)-�S���O�a��FB���zŀ�ǵ��*� �i��u�*��~ �斧������PѨcfB��b<�^"jU���ǚ��\���f&j5,G����F�S�T�t�>s�6��"�}��}"h�_��G��Y6r�Ȧ?Z�i����,����R䜣_�Ǆ�э�O8�D�	�?�l�%�� 4�jR	���P����:� ���j-�p� ���;��}�Rq��]�:�������V�-����UtM�v��n_�V�o���r�T�1�Uŕ�"=�򧦹�9��e0��w�_���r=9��'NY�P�!~��Ab
��\e��=]뚛�]�?״��z�wt� ���tT���C&k`�#vQ��h�" Mh�����[��lF{3��eI��WF�EA�5>れpaHD��]�B�`td"5��*B(pkh�<�B~j�����k��i�M'����ü�P���?$s+)[���a�p�l�+�ϙ�L4!����yh� �QP���tX��*x$�b�_Ɨ���c�x���D��3�Rف_s�A5C�T��J�,�{��R ���^�tg���*S���U7�FBpT�>��UC�Q���%��k��;��j3n@0��4�(�Ӽ����I�E����(b'炽�܀T(q�w�9(C�[�6g��R�}���B;��-jUڱ�������֬J�Ʃ�)\Jb0���l��q���`������P`E��_|v2n�wx\Ġ�K	���]r��Y2%$���/��~2�wG��M�픐E/JH�����C��q�ޛ�$t0��������X�<z�8����{3�����
~j�8��Ѿr��V�����f��mC*3��&yj�G�����w�M)�Q:��%����ŗ���,���{"R#m�Ĺ�&��7�A֐%sۏ�~~eG$45�K�vWY��P�)@U������OP{���	��e�w��pr#� ky�_ީ��H�uT<*FG��I�d����Z�W�noW�z�QB�g�>���qÖis�f��@���D��Cl������k4�I}�z���*�K���[	�I_��bz���.�BT{�����j�8��P�_���V�K/&�NRTQ\��S��qf�:�ш{��5�)V�Ή��<�m�#�F���.yn�;���ZP�OzF��S<�:g3U���p�o���,��x�e�C�nüx��h�c,oM�V���2�1�I�����hs��
�{�>Q�uB���E�t��uq�����ک_�J����)w*�y����⛵��o�#�����s�PBu�/�i:�� q6����O�����NP�te�\(�k2p�am7�Ty��ű��Ii[���7����J��D�+e��|�Z\�-0cdC�Fw�2qD�e��"�(@��?U/�\�(WCO=�p{n�,���=���,�|�����C~�J�0j�m�'����	�0�z	36FO��3�R�}�H�@��Vh+��ӾMƅ�i��{W�����ri���|���b�b|�ǽ�I�G��6�̤�v��2z�V��$p1�@�N�e4hS��4:8��'�g|�E�0��E/�x��'#�}��R�5�E	\xhiVT�;��T�E[�?w��C��=I�FsM��)�́i����̀�w�LT��7�7���b��U�8�jw$w���s"6&߯�����'�؜Mt�ʩ�.����iJ�vө�Kkʄ�v�us�0��;���J�O=ו'sxȆ�Gx��S�J����P�#��_�����4!^�T�i����Ț�L5.]�����F�.��J�K
b�|$ɜ�c����Q��u�K,��ز�r��<E�|e:S��M1��ޑ9�ױ�e؎���zDM���Q�.���Vi�=pҿSA���}��؋��8�{_&%G9 H[�j��^M|F��c5�Ϲ
4)P�0"�	�-���:@_�In W� +��}�<�/���	W�ۢ��i�