��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����>�S��fI#�l7x%���$or�#�6�y���N�i� �D��f(�:eǊ�` ��S���^�mBƱYjA���v�0��kh������#�v�(#W��ux��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf^��$�i�g�Wɐ�)
�Ql�Y�+6�iѰ�^���d�u�.�Ye�ZG�$*�f�pM��Y���f<���YB�H6]��^�8�G{��:RjeQ��2
�ƣː��5JLO%/.�)����\�
,��YIw_�aJ�/��]b<Q�	��E���i��U=wx�-Fe}Z2c��~��=' ��j�z���Ҫ�dC��U���=��/ɳ��^�+^ ?� eZ���[WF�ד�������a�{����A�����t�	s�n��~h�iP
�������P�iz����d�v�W��Nn#yx_� �Xh�����w`�`�#ו�=�9y�U�B3���k����[��_G����K�����%5���U��;��v��������p${"`�$����?*��6���#�6I���jѻ�:��C������O<�-{5�̫�$�Ɓ���>A��J��k6gr>fR�KA�#��~R,al(����Ћw�9z�>��c���Mr�ɛMR����|3o��ב$�Y"�Wھ'l�T�l��P��5nP���+�ł���M �KY�� �C���r�QT�+�ʻ[.v{��8�f�?]�K
�,���c3-��^�Y�Z��F�3Q�>w�S�ȸG�?��$�?�[����Qئ�kd+8:>�-M����͈�ꯈP���p��E	Xt�x�b1x1�!u���k(S't�T�bA�a����SoGg�
[�	��cP��\�}}����O�6w������y������MzEWS����-|}L�<S�ߐۛ5�:��@z�����������t[P͘��`<�����>xc��+.�V0����&4:�����r����0�R�u�N0d���K�9�LhÔ�ب`E�������iW$�mt���u��՘��\�r!���7m�XL-�d����2�W����(ڬ���D=}��[�X�M]�5 �o�ĭ�OElAX1-�f/(5�[�q������+ǎ�|DQj8^6w`��q�Q��?]c/���ĨQ�wO���a�Y��}��ܫ"�{cS���!�n'~�;	�I����C�||�'��g� J�WqBB"�Y�������l
teΡ�F���B���0�d��ԯ���K�-�u!�=g�t��s��Aݐc��Ǧ�;��;Ƣ�+P}%NW��;r�Z�Q�	��l�DI�M=����/�7m5�"C�h��Pc��ݾ�m����F��M��U�1.����Lģ!?;NQ@����Z�\���i��j1}��y���;|�u����ix�)[֒�{�;���xa[9,i�NBF�`�f@l�I�xR�Y	�1J_�Ӏ9��cw(���tf%�
Eo��.��0����^��0=a��Ga z0�(	����nű=�*z|�Fl � ��{%�|�R������@�F8��0.�=Z�@z-m a�p:� ��E�i�;g1��"�)>���!F��>�|���h�p�֚ȵlo-8�������4���g�g�4>{b*]U�]������=�4��7�-���MV�"����!#*�	��Y#F�V�ucʞ�E�0]M�p�7�ي���y<YM���Meh�!\#��O�;Qk6LtCuc�9N�o�Y�ڒ���C���u/�&�)L�Y��+�6��^�^=�"3�����%q3⹹�Ɠ�?�$��Q~ ���r+�i�{�"!�ڪ�7�=s?jt���S�)U[����ucS�������P/�@�7��YoҀY��`;���	����dϲ
98Cg�+BK/����䞤�Vjhl<�l^�#e�DR���3�+���+}��+���X�Q�^��0���:�~!Hs���x)���l�n�.֍��E�H��)��9vJ8ߋ����� : m��6n��4���7��ߋXm��H1�ܗb���m�}���5�c:H$J�a��U�����>RԨp	��(���0�F����|姹����GQ�������P\D�7���s�5ޚb!�l;(���n��"w�kU��6;�%{��0]$pk]��C��އ}�5K���s&�Sie��`e�����i�?� d�}�s�h��
�M|j��m�b`S�~�	�p����7���IXw��	H�n|9�j}��pȎ���x+��A��XAx�ʾ�6�ߝ��;��|֡� �+�^.E0H���.����zJZ��X���|�ɯ,�1�E	g(|�1��̓���am��5����c�� S�?Q���ݷ���1K~�\�Mv�0`�Bw�\D���j�5cgYƸ���.6�2��Yr޴�-��w����\ �����U�FY5/�יg������5�����o���O��`�ӤO/7ȣ6l�a@��������P�Gw �������w�ت��e��+a�B��E�m���6����n�~���W��-��E��Z_�	�we����9Y�+*@��c��|ot�ۖ��5a�cvrf q8VvJ6Ė;so�Y�F�̐i)�Tz��&!I� �=�H����n��CB��ć�ɏt@%��1�g�3Z�ԙ�@�/�`>Iq{��d],� 9��l�?���_m̳j�do�fe.D�n�s��o�]��/g�t�������F5$$��,�����9y�q.X����5�óN�����/�"/U���>����[1J��64<}������~��\�+�e1f�>��>�~�J�~a�vq���e�x�n(A-����rU�qNa��E�����#���Pw�(��w�OK�h�7�L�h%�|�K<[��r���`%�9t�!Gʳ�Ǖ]!��-
�-`Aм�~��܍���J�x:\�!3K��#v)c&�_�����;��v�,�����l� �bPl�ю�Q*p�N�-vqoGnQ��422�8 z�.� �j�[�V�=�<7�)j�+�R���Qm����O�PX�GҖ������(Z�K��MQ��KZ�r�z���@�����5 ���2&�P�;�o�}~%���ǝ�<7�W�K�?Q�/�I�ShAϬ�iц$0w]˯�C<L�`��w��~sIz� qR��!7�Y|���V��Nd@�B��H������&f^��.��.iy��{z�?���_����qf�7�����[�_B��������m��?��M��G:涆j��p`X2|;#��la^z1�o��Xm���i�B@�ˬ��|���2f�).Ē�� �!P��_�����6K��Nʴ���IQ�)xM��[�z���������#��x�2�B���v�ᚨ�|8����'��p�mu�}"J���<���8{�G��xy~���d�j�B��'�S	���!`6�'��q�q�ޓeڋ.�}��0!��H��|�ڕg��> |���o�vs���@&�b7����.���M�F"<LE>w���-Ӣ�'2�z�!3�a�G��%�U>�Ht7�M!.n:>��կ>/L �W���I��s
Uʬs��.f���ܥ��&�%�=�H'�~ᶿ��,w-�<��_�is��A��=�`��Зع����|��Ny19A��U�m$��.u-N�a<ß��-���p
��9�OQs���pF�D��Z���
owq���JK��
	����x=X����b\�|2Lo��<��$���d���vT��ڭsP�Q�ux��.(P�lSW1��f�����F��ATL>�X���;n=F�
��r����÷���6��E���d/�t<�N����R�T�J�����q@��l�T��xk?}"R���`�R�f�<�<�pw��8��a����~Wst�j�/�kڌ��������Z]w�n6;���L�l���`f^Z��ȰF��M�fga0Z=��Z ����ʎ� �7���3-��Û��7����3��ܮe�k#s�@����6�� �T���Q\�a(��#������9�C�����`i��_|�7zi{F���U=��CΓI͎�2GtT�?�e0*։�й4!���_�&�ۀDRɾC{}|�Qz��j�c��Y`L���?���ѷ5<>u�>�ވ[G̰��<Y ���xqߓ��I疍�e��ӂ��*��h��xLF��-���
�"	0��%��6C�j�L���?2��`]#�ء�-/���J���v�bz����ҷ�� /Q5n�	���Y�����D�^_<��� �����Ck�(wP���B�"=ˏ�
؝�q���@O��0�ә��o�Zܐv�F�M?���2���zc�@�A�f�v��7���.��o�6i�!Vs^t�l�A}�m}2�,;�΁���!2�3����(�=g0��a�9H&s�*$j��}�u:)@�e��޲����(M����:[�	����U�
�\���6y�^����+!
P�����N�������[�-⹏V����o/Z@��Ƅ��=��U�OYߎʂ�2a .��4��
���A�#I�a�`�5GJ�,���C5�	 õ8MT.�8� ��.Q�&����*��8S�K:4�(*So��f;o����g�+�\���腔w���W<��N��v���k:E��2+�H ��m����M��4a�e>���B��c=2�2�s�'��Y�,�D�f}�\#����G�ܩδ�ˬ#�	�߲���	P @(R;��3�p���>G����[[ס�^�hl��fXLw�BGX8��Op�A��o�7@���F�'���tݖ��A=.�)�CQ]%81���V��h �
�)�ɤ���9�ybR��޹��̣�~s�����7F&�@��̉�����ZX�����:����KT�H���A��3 5%\�D�.���b��e.����@��9_��6琻̧����b��U��|�I'7|�]I�W�;����j�hV��B���`F"`�Jxl��I�2��l:����'�L'�)��w��b�G�@>��VV7���gE�'V���<y�g'�TE���a���ّ���wb�-���BLr�]B�`J����5�iW* ���W�lV� S�}�]Yni���7{1�ށ�y��iJi�/F������*/5��P��%�ݐ����Àu��N�H�4�pY0[+)@\$�7��s��᙮��[���@�߸IŚS��g ��6�ivt��ҧ:��Ce�")�f��\rXt�'��p��1�!������ܠ�ï�Ġ�X����$j�:;�d�t���G>��E�8���R�0����%R=�� ���")��`S�f�
L�N.TRDþ�НK�i�f�
��mɃ�u��|7���m�̅&�oI�$�7ǹ+[�!�.��Q1�3M��p9z���u�ˌL���nqK`�ʼJt�[Є`4�<uH���,�%�Z5�2�1�|�#������~@ �:"ZrW��&XP�F{8��-9�r{y��R־H@�c���q33�y�6�/t��(/)���(���ы�o�������fl�{�aj< ��C9�����%b���i�Ɯ��&��]���r��1|�w���l�0��2�7N��N���e������B(+h�� �c��?}+N�jĄ60�2��{ˉ�������IJ�,�0����]k�F���1]��o�0���������5��#����VK�E*�U�>����S�7um��t�X��W��h9K���m�D�k�����<���.5'o(�|�j	\�QNw.Ws|�2�5R��
�����V���dP��H�FL�6`ޚ�u� �-9p���V�U��q�K��A�ʢufpf�{��+��f>V�p`�Qz���۳Z���ˆ�[%$�m�4a��%d��S��h�U����uR�ݣB0*�\O�Q*��R�r��iHA�T�l���؄h�M�O䀮f~_�p�WE�c�Y{�=�g6.�^Ku�1��nԐ��r��H�����7i��ׂ��/_�33,����l��E�����p�4��`Z���Z�F�I65M���z� x)�C��,LQG9X/�?y��0M�ѣA�)����ġ�����	YOk�o�m��\#.	��]w�� ����:��bP3�O}x8hQr@�샥�������.<�1��<G�p�W���
�=�<e]� �^�P��z���Oד�?�nSm`Z��b0���;+�u��J��ߝ����ԛ�x�β��%+�ܕ��|b\��u��"�����j\����� �R���G%�FNP3l%�72[7wĭBcr�5�<e�:�v��2l'+��a���ny����S��J���9���-���l���p� u � I����ك�; �����6@!	�{�/X��АN!�^�?F��P�y��u�\��#�\ؘ���衊B��(x���n����f�Mڭl�8�p��5�8ʤ�t�evs�S�f$��T���]�>�Xd�۠�F���(��v4�J�ĳj��>���8�>H�h��8%�W�41�����HJ�6�Oi7N�/`�~��10��t�K��i�U�0cI�0/B2�,��*�e��k�9����]�wd��]����8HBܴ%���q�}Qr	��͗���?i[n�DL	/�d���|4���t��� X�N����HG]�P�	bzdq�,��<�\��P�T8��hm%j*A�G����¢..�SC�u��ք��E�V��g�*�1�h(�C�;W�,yE܄�9�*�8@b��Ӓ��6��oQQTCk��$CW|�߸x��"1,�O�o��LqRsˍy�	zI�-�~k��	�"�%�����OT>yx�=�~�5
��e��Ox��B�������H�{;�0&7��j���	��Y����K��/�N}�|�S��:���>��[
 >=~Ozߒc��o�D��Zpl�P��0w�<�m���?X,+��ű&�60QN�'�E���F���Y?�T�
�%�@��v��6��09�J�o�lr��2��3��kͨ�L6��|nd9xC��%�,X���Ǻ?h�����ㄫ�7�ދg��`=_�~�l�._��V��^��o�y�]q{cE��Roҝxˊ����9�ݫC�S�0���� ��?�IMAYfvK9�6-*F�����?����L9�@2����y��&L]���/�EԢ���>t�3��Fa�9���[��+�ᥲ6�p�g��[��^Mk˔�{;��;��=�mbw+��̜�R�:�j��%�d�2A��L<z�'��K�����4.o��ÓɅ��}��(Ύb?T:�-�ĶI����ʭ��Q�9Tâ��l�+؞,��5I�:B�&@�8��}����=�1�Y7-�
�+�(`�0�'��l�ڽ�����)�:_.�s�^<���Ѫ�*5�8����<
Gw�yc�a�ι����n��1r���B����������^i�b�/�G�o�TE�=2���f�n��~Q�B'5��z)�������Q$<AP�4���֯� �'�li�zQt��Z�ex-�x��ADkx�NL�A!��ȟ�KA�|�)1U�#�h�_�5{��H^ *X���Ӂ72��3w��<X�xf���������R�e�DQ}�8�\��^�}���\����^��6'�U�n����fLAt)t8�	
l�gfs]x�dc�i@oGar@���c6�k"� �&�	) R�[m��2�A��k�Wzŷ�&�9�x��Z2o�n�Ô1gʟzG|NP�p^���_4 k�N��%/>�y�@�6�\������.S~�=^B``�A$�&*������E<-x�v"�V���V�P�ʲ�@T��^��I�܀�PEn�՛]J��t��߱G)�uY�&�i���<��w��r�2��FJ�9{
f�L/�������\�t�3���\��_�vѫ�^��l��/��.�O]�0m"I�&W�kNA��˪�����v��nϜQ�������	<��(��۩#a�.+ṬQV�:���V�HR"�J�=��.:���Ȝ>��[��T�E��9�I>w�%��JN�	V���dYj,���&2���1�c?Ԟ\zK/��tyvH~=�#��ڟ�rk �Dr�K�c��������̓�T����;2�����ǰ�Li����HW����*!���ߐ�ûsI]��� :E#I!��h�l��B����%�z����(g�#�㣍%f���&�˒�~���R[�Y���]��_����s�(�r������.8�?šC�ߦF֫W?�?p�b}{�+��{�n�YDH5�K4��R�eLp|���kNsNW�& x�pT���H��vF��pZ�F�o��J��G��*��%eK/�W��R����<tA��*o�i�U�� ���]� �V]ɰ��t��ȚA58*��V=��eiWZ)��"u�c%4/����G��ň�M�9q�:u^�p��ot��0�tj6�v0��y�������48�ވę�f�$���A��3�@��	ԖJ�sQ����qk>sg��2�!mq�G�_�2� V�-�b��D�6G�/o��!��Y�\g����%���	��w���|2}j�~5?^C�����X���UX�en] ��Ve��V¹�I�ڣ6�r1��ӵ9�i'Z(�I�W���*;�N����k8N˭=�j��}�3�5�Ys��ޜ�}��#T�y�C�3�v�ȱ!w��j>u��q�\ģ:��N=�C��cB$	?#HoY6����{h�A,]#q�㒔Y���8 �+�{ 3�O��:|Y+��r&�	VZ,R)���v��L����]�D�ߕB�E��"E[���V��HdK8��]�L�Ԑ��7�������y������	X�.����*~#�gs�w9S�Ƣ�Ƅ��Bj[%��}�}Ic}����JF�FF�:�S��հw y���*�LT{R���Y"R���
�m��q�A�_̮���! gi'����H��2\�6G���	�G�L��.ՠy���]=��:1�@7s�itn/���e-�ht�:��ף8�����[C���Ls���5	7K��Z���u�m�A���B)G�&#��LyI7M��5�z��19|U�Sp�GeL�<\8ot�8��_�~�;���u8�)��UjY�L&�[��L��Q�.�A~�)��\H%(�ea��mw��?ΗQ�����+?�6�h��a��W�>SWaJ5#0�y�C�Fp�XC�u��������3�?+��m.�za�.��gb�rƅ��T:q��ҿ����y%��g� X"� ϳ�r�e.o�t'��|7�����H"����<]ŋΦd8. T�#cZ\p��S�eq*�bBYHX����'�M|�M�>oi[��H��+��2OZ�*�l���	Y����#�(�����;D�p`����k<*��o`W`{�HKc�{�`cG^���]��.�6Q���hb��y�{.{]�#Ŀ��+�][=]�M��4t�`�Di�S4����8֢d;gv���ex��?m�[��� ��g��'
�ՌP3a��H���<C�OCS<���rt ��m�M��i�I�/ב���ha,,d�W��27_�>�3?�ʀ�Z�m�:@�ԏ�?T�{��?^�fг��7����
�Q��f����0��%��B�W������Tт$��%9��+O�?�Wv~�cY�����I$�0:
#=��P�V�]Ү�^��n&��2v8�C`�_���*��r���}A�5��f��5eU��c�4n�>���Pқ���Զ���W��;$�X�
 ��n�]vIb#Zg@��Ysq>�48�L�«3��b�6%5���ԸV�jm�)���f�iT;w���Q?��Y����5ٔR�S�#@ި>�e��� �y+��PL�,4���pn �"2�7(�-�l:V�&��:���x�r����1=�W1q
�.!"�{���x��=�z`�q�Ω�9����m�")4X[!�F�Slg$����1?��bPۄ�H�Hf���Az FZ��4��s����B���ѣ˘2�Dh�b�{[$tn͜�t�{|�Bͣ u���{FW��	�bO�h����^aaèk����, ��e�
���>2�0�jc�ޭ�ԢƅsP��� u`�B�J����/~.�Z(��qG0�R��D!O?�<Cj:MQ�=!JZ����*x�1�	]�Ig"o���4�T�Z�4���<@$��pmm�61�uf\Ձ��KU}��ke!�PD������#<r�7&,L�M�������s!�t��79�s�攝0�bX��k*������E oWݘ	�s�d&☯_��suy�TY:�`��������׼��S�r�.3��������j�FZ�,�ȅ�BgòY9' �~$<kz��}����g^�{hA�.�.ف{�*�"�Jp�N2�{������B��c���t�d�Sj��;�w��8����^�GZ)
�gA�#̞�ЃNΌT4���!R;����h�ё�PJ���E�����eo���Kj���*�MLn�8TK᝚�j���,k
�ݰ�a��H{�zv��5$�ZQy���kR(����|so�P;b�B��4�T�%_Ƙ���)�)���@��-ax㟚͘�ya-ԩs�zRa�����ڞV��cR�:������,�H��{R�Fޖ $�m�.x�ҏ�Gh�Ǌ�!v�8Pb�"��	�r�I�6A�p 	c]�����T[<ȁ��E6�Y4��Q`f�Ļ�.�iLufu�����#R`v˕V���e�t��\���Q���[�ڂ"���$-RI�n���X�9|���õ��e����d�QWZ��c}vwu�h�8Q�>ysOV��,]s�kr2)��8�@���:���׶�rS0�*�V3�)��>�F�Q�s,ɐ$8�b����/'��Wwx�f:5�.��@�2�����R=XY�z��i����l�GLۂW6�v6�NTf���$)��Z�%\벗�z���-T�:aW��cEԖ���R�Gq��0�nc_v��J\w����Ֆ��ai��˰�#�LG��D���!�t���!���`IP�e�hW��z9�	 �
�Eq�U�[ǌ����.�(�aݬM1��U^k�VO�]Ԍ�d��#�I�r3�&��M6�z�}a����	J�F�{7F��1e���鈃��c����eH3���칆x�*��b
��φ ��	+xC�]�M��򃊕Ii��A�pE��}�P�6{nٻб�@J�������T�o�����	��|y���/��	S�q(Dߞrh2O�w�	ES�-�U�+�����䇺��Xn��R'&I�ӛm�P���H�	�Q�vŊ��èT��iE!�Z�)p��,u����a�ܸ\�UX�{��<J�j�R�S	���V�}g�@�����dٱSz����_����Ǵ������K#������=���4�^*
����1A���_i�����!�(�7�KY���L�ܩ����0f%xv�$S("��&��$��&xֈW�o����O)�G9�O$�4�ZU|�*�����J�J��=�r��Ds��da�ޠ3 	u\�c�~�qv�R�L.�!n&	����[�퇄����sx�o��^�	�|���ob�]��z%��=�OvK�]�y�R~QElg�z%��"٬) ��j"�Lh�*��z�\Q�K�qή����xc�D~Ud^F�WDMXb:���K�=B��#�Q`WXà�J�n�0cYlo�=x$��6-Je�����	��ak,�Ev�:�"���t�I�d(:�R�Ck���O@����ȍ.�G���Z&7�7U`_�HA�C8oԎX��Җ2�ى���g/r�t��2�:���	�tJ�P�j��}�d��W{9�ۼ{M�g#C���k�����{�Z��υm8^���9�T�6�d��mc+gE���p0)��!T;%3Ҁ�"��Z�w"����[3 �0�[��(���_�	���״�ݨm�������V�7ؖh:���&���ˆiq;U��o��g�:��:��b�w���c ��bBD�B�:%I��o�:�T�g��;��tW�D���_�_�rZ�͓/���ٷ�!6]�tN�gXӨ|�;(ZsPЬ�
�^��[C2�@�z�b��R1R��#����]VXZ�f���`^��k
~�V��Z2��T���d������ix^V덋�Vđ���+�?�x���u��;W^`2=*k��bs���}�'��бf�8�q����N���8���3?�ˊ���;;�����7Xn�� ��
�Ez�kϲ��`�� 3S׿�:&��`}�+�2�+�����֟��qJ3F�iF�g����S�kJ���{�1n��I�g&��7p�\������Q� A�^@- ʓ<;�:P�B�;m*�~���#ɇ��/�y,i!���DCc�/��T�������N1=��dflhy���{�ͤ���;}���vL.�Ys�d?-��k���\k�P��?�_�C$���D�%��I�@ H��0W
,�ڠ
E3=��8\�T��݃p�;����������(9��� v��U6��N�CgP��%��҇�1:PT$삁WTL����D���<K��W�
�dRѿ�B��ؖ+ש��k�tCC~�5N�÷	�b�
,z°��Ƽ�f�ch:�;'�m�����!���� !ڜ���pzB7�
���w�khdq|$x��v�|��.W�SRf�Km�5�R����f���z��ida߃���k2�~������z�F�}�G�ɝ�ط?����I�{�gNߚcl	H���Rf���XQQ' PIR�����S ���e��l�ѥ\�3e �,X]�o�?J����/�=l�f2)�)�M�ŭ�Q�"9D�����[������=��;=R��*e��3AɁY�C�Ï�vS��N�+^�a�9�	E|�w^f�����M��KCOK�N��8@zȖӉ�.,�޻iB����YMT��aM�C�(i��Dڏ�{;�{U���j�S#+�x(��o/������>WU�q%�I}���Y��m��Q�
����[=$�ׇ�x,l�v��u_�2�p j~�W��nv/�G���uK[���Jmv t�a6��6~�ZP�b;�;��K��ّ��r�yzA6h���P�:�z��
l�� T/�C̬8tU�8��8�&��Fkkp!��2X��T�{���:�]1=:u�}n8.�1�n~���\�Q�((K��u-ոN����(��Glއ��8�8wLJ|�D�^i�Ф'B$��w���&ǝ.gK�_���у��p�O8�1�=љXM�m�	b����A�]}t,��+��ǚ~XqDGpY�A����rɤ4��١Ҝ7�p�����Jn�J�r4yW5Xkӎ3آ6����Clw���\�v��<�l��d=S����}> �#H�-ƣS"n���t�.Y�%RS ��}6�t��#�� g8<�L�o����1��s���WdJ>�&��\�޿��\}u���R���B�H߆^���0O]���l�َ��"���s6�ܣ�k�� �t�*�3�s��)������q8p����{)�~^آ���]#��a%�Mo���Y�Ky�cN�k�^d�4Ru;*5��K~b2�-	�/�^5��Zz���
�f̶��ͤ��6�ߋq+TKs����5T�#�:�ݻa����Nĉ�"W�Y��9҃⁖�E0!�Bl�הe/wb�Ow�;[�g]���!�����]�=���E�k3��!b�����H�KZ7���g�p�ju�D��r��p��ﯛ�[z!р��K�wHi9�(��N����s�s	n�Sc�;��a�R7�_xf���V]i2@?W<����h��M;=۶D�(E�NAe��a��{�t%� 0�����X�I��P_Z��&��>!����%�<P�y!y�9��N���t��L�y������M�J�:3�+k׵�r�
��q�%Z�d��lW�ۗ�����W�a�~��b	��5�=�;~���������RZ��o3���;\�����ï�3]����]��FL��m��ק�$��7X�%�������6Jk##p��]s_y"Zfm1\�p�d �r&��� D�O��ĐMll�
��:��z�S��Y���:�r�:�)yF%�м5�$Ԍ��I:3B��l���.���	�O�#1�H�Д0��" W��R���۝S�ב�	,5��F�n� �������i*F2#i���ܽGo�]�����x#[n����d�Ӊ��H"��X�����	F��L��<���i~��ޜj�kɵ�i���{���V=\��y���
��Z7�tj@�������7B�D/dǷ�w$��%���פ(RQ��nu�] j�p��W�as�'�6���u �L��_r �� t#.�vT��mF����x���<� F���2�58�T�YďU�q�:J��陂H��&�g�H��9��7+P]�Ze�A1�#�̿bI%�gWs�d*ۚ����%�P�� �������	�c6�9��p�<�w��N�����ș������Է_kGϼ6S�������O׆��'����vm`�;@�n@Y���˪G�v1�C�����Lb���=U��#y������{K��r�r�d�4O��E�'s���	�v�
�]��H;j��TN�"^�[/��C��'LŨ2�R�-��{��e��C㕚鮷E�`Z6:jJ��rr�����}��2Brr%�o�C��ԃǲ���b�|R:˶�c�*�M�'g�/r�'Ʃ�]�!7A>p���;0�/ꑔ-y�ksY�1��F��7��/�"m1��!���<��,�N����/�\��:�\xx����[ˍ=g��t\5���~����F(�4J�E�/���皞��	}rk��p��h�g9B6F�9�@l���A�Rgђ����VA�	�L������ 'Ju{��x���wq�я����ў0���!�][��beҢK��a��7��e/�.Fd޳>���_:YG�i��L��j�?Qu�K�L�)Y=�����z���3�"=���.ț^�0��J*��h�F�ĶuU��/�kϧQ�y���9�!��ߙ(�l�믨)�>͵�޿�5l�D��w�<��p��5?�k:�
o��2U�,�IҿH�@|F��v��։��ŝtM�.�`$��'���Oc�^�X�M�9[h"�9C� ��b[�E���-�T�n�8M��:����F1�k����X\E���dTP��%ʅ_�5�䋌�/�����ț��)�+)�x�$���ؗ冫�n��ʙu�d�>٩#B�LT1{z�Up�mbW�M�@}�Vz�9���\!<�H�*ӵ �v�n������4G�~���ָF����*�e�dhY��b�}f&d��J�knG F������3�zšv���u����3�0:�\��MB:[)V��)����:�:p��"!y��K��HD�ko� *��,e��\>�N�W���a�S[�=c)��d7�}��,�f*na�U�Ϡ�������%�����x�!���J�$�Є a�x���D��J ���1ٱh	�67���Vҗ5��%C�pi��LdRcND� ����N�1��>�����F�hH���cW/��/�م��yĲ>L��8󑵊~�ፑ�����i��	@�]k�3�(���c�뽕^���3�^�A��KD�!M�e��2��T�koOGvU�(���F��	W���0Y���cd�^0lW%���gX��@l�p�1�m����d'���#lJnI2x�r����N�O���^����&��K؞�o�Vi���\�ƣO2f[X�I����<�!n��sK���/8�[,��]B�㟉���,_?	z���?a����^������R��
�,r;��r/6s�}�����(�c��Z	'e
/4���VFb�Y�����P�:A��y@Y�� �4/���v��zb�C�U�O�s�����9�V4&�j+[(�x�c�\�@�o�)N���]��	��Jgc�02��mܿ��@ބ���ȡ��x���[R@7��_�*N����f����K���V#�b�v23�a�*|���E�2����j͙���|��d2*��;̝6���6,	u�e�W=�;�Q�f���1����
��$
���)s�=�7_&7�W�&�����?^�	�ݦ�)��vBy|}8)��fT%��q�$Ǫ�_�DϘD��'=��ϔ�����:(/)���/{3=4͌m����J�$���Ԙ�d27�B������4��k��?��z�^����P�(��>6�}�*����[?y7�!cgD���K��w��nD+K���/@05i��w#nBN�:�X�?BW�Y�����.�7�#��w�I�'C:��
z�ȫ��:������AO�Bz�Ğm��x��^������ �9����!Taír���T�f�D*��z�H�����j�6M��)
��Q�'|��� �3�\ex0��=f��l˄�%�n�U�1� �Z}~ �J^j��wd�L��S���5��"UwU6"���vO�0̜ܙ��kc�� Z6�x��K�M.��__�/�p��"N.��������U7�{��P����8O��k�!�$4���?�Й���v��h��v�~Is�{iH��y��M��⃴�V������t�)Us�(C!�Gqm%�'q��9k�+�a�^��Wdr)"רF�*�{ �y��g����Z�li�h8�r��3��$�r/]������c�k���&�yu���@P�wy�1YI��[G����_�4�xFͿ��}�v���x����xD��=:L�B>㞫���@�IE
�#[�v�E�b�1H�B�:�����p��h0ut�1нg		�w&s$�h����<.�ߍM��j�@x�P ۜ��v�r��o��)�Ȥ�0:<�}��Զ䠔�db�Fퟓ\^�1�Sw�_��SA>B!�P�:�?ġ��g�	��qo���[�1F=�Sj�L��N#8[���6JC�=�g3`W��LܔFggC��S�w��dG��k/YӼ�7q2��)�0\TM�ho�v�*�gw :Y�h���u��Vy$Uw��k��F���f��PbΤ8�d�<;�[]"�m���'�h#x�sC<��9'����' �mCݞqr� ��ɂ���~x o��ise[�J�H�S��f,��*��D	��:%8H���@��ͭF���s��;d�/����5�0ē5���Em�غ��y��!��U���Ł����|��M��Fi*������Pd��=�W��;r�"'�@`�vD۳�_�<�B@&װ��e�Zה�(H���dt����E��s�?!��B8i��}۰7�C�N���z�a���y.9�A���)@�ü{��A����P�i�B�3VZ��~�{�j�[��ĺ)ν��fM>�Bd���~�A��d�N�R],s��N�i�T���h$�TJ�c_���M�2�j���Z�͌�)A�q���\:�Y(u���QŗAX ��v=պ�#���Wtd�*4��(�;����~!}�<�@�/���.-���3$��)�h�4z�^I�)����S��j���&dz�֟���ٷ9����rE�d�6w6���	٭�}N '!F�����^�L8r#x+��m�Ҝ�J����d����֟K��Zn������$Q:�������!y_��HP�.�B5�M,\�p,���^%B�WI����w(�]8H	��ק�=�#��ج�u��0gxq��rn�Vw3�*y�"̮������X��D\ur�A&��T���⻠@�O�}�����ߘ @ �`��$=�^�s����˽r��Z2^sxI����<WP}\�r�t#�.�Z�Ԭ�̽T|�_L��:�A�ӵ�eϧ	���v1A<��,>�k>p�[�����!5�-��Z��T�qL>c��-1A[n�u�az�� �����x�F��|�L�٬���G��LҾRg��k�N�£��̠�*�|^���1d�`w4�Dw#E��aT�B�����j0OШ�B���R辅XK��b�9�Vd��օO]��a4/
gY���p��Dʑ��B������}t�H�K�Dt��׷�'~N�k���(
q���8�s�F�j�lB�m�|x�#t����RWP�E$`�8�W�r7���ӵ?-gH���M�ȺO�*%�f�b�m�[�i =O��j^��"��"W�4�)���j�z *�a�~#Fn��%Frg����z0o�ck��y�&��- �.��wx� �#4�\-�a"e�iq�V�::��B1L�a�@��H��#�<��9��2hY��skL���uex��sǯmOO$V�9�N�Ms��;{:6B6���h<A�?Q�%��i�(��|i�~9��]29[������e����P�5�
K��ҕϐN&�罏�k��J�MϦ(o��tԭd����m�N�r�}��z��a��M�Y���R�D؀S�
s*B���o�!��0F�Ш>�ʿ��V#���HG�E�맒R��[^cF�5^���~��y7%"N
f�"���	�}��s� ����r��IO�H$�,4�-�#��¶x�(�[,W����~*^G��ޕ��/�G?��8`}��R�yoz���%�r��������^_M����8�m��m���Q�Fl��	����6��P���"��ܐb��v���
��\L��!ڍ�//�A�؄pxxLV��	����w��/�8�s\C�3�-|��&����j�UK������e��E9RRr�ia/7�tI�%��VX�{������WƤ�Z^ٲ_8r&����F^w�&t��(��:L��9H~\�+��-Li�
�	��5��@2].��ؾ]"�2~_GG��Q����B'da�����)iֺ)iSL����;��-k�9}}�"��ɣ�-�k�p��Qg�al�0m���`�̩��r�����ᵕ��F�D�inQڰ6�@'9M���>�5���+O�b��ı���]� F��fT�z��i���\�l"�q0uB�q�e�,L�@ְu �"5���hD���E��m�����]�)L��`��{(e@�C����X\�p�?�̟X��@�"�C[0�����S�KW���B����Y�qTX"`=�����E87��	�`��4qW�ϥ��Wī0�>�"�(����3�eh� �/���P�q�&��*
UW�a_��F[|㦭��M���j��4��XO6muv6�5�vX�y���V)��Q��P�e{���u0�x��ly],���ܜ������!g�~�/��i��p�]:P/a�f���P{�B[KkK�C
6�,�Ʒ����D|}h�)��T����3�_���+L��,ӣt�2Zj����N��k��$8мQ���[�����_+c>���=�
��J�������5�B�Z�l�Ա�|��^��>�y�-�\����6�;�yG�ꞔ��m:��j�(;/�<��s-J��Ҳ(�v;��T
���=�`�v����@���p������й~��*�e\u�X�U_T��#�/5dT�N� ����*'�?�`�?[_�9�*���۹��&Q��fA\{!�7�m¶ʻ��r0,�,� �J�#�0��|��n�cB�UUa��lB9�-�������sy#���r���zw�@���r�?���/J�]�6�#��Zws�I�>�_	���^T3"q�˘�
$�;Z	����4f�I��rڡM���<�� =�!@l�'����t���)�6�����sEՒ�̩V1ƾD�J�X���e*%j�2���B�ZQ�D�\�.��fFG�Us�)stS�ϰw��4�cu�g���0�� t���!����c��f(*����k��g|�	h�7s�q�PMuԄT�"�+�+�+X&��K��� ��rmpR��3Z����v��P"�O8��a=��6��:���$@x<� ����;�KJ�] g���Ӵ�!��������]O�Q�vM���	(�9M*��i����ƴ���*a����a�X�1��@�Uj/�����۔f&-��)js�m�3�{�r�9v�	`�~��{�m�J/Nm,�\�/5)�r��F�}����o�lo#�^-�W���Y?а�@[��K3)��HH��6O~Z*оy:��F蓊��g�Kh�<K��
�����Όw�r�,�fv|�G[��$Qq�~�#�^����Bm�5�~�F���P�[�qŎT��V�{cBa�EX���äu�#�q�;�9�hQ��뫛 8oM	�����"�y��$>��$,�2@>I����"i�K���p��?�U;/���^5t�Ĉ�NLtN�-nс���fK�oq�TݭȌ��LR�i�.��F0v��la	�@�Y@�MR��X.2r(�\g�Z��Ͼx�Q���ǥz���w���
mފ{�b�
���鈥eP�穻z �(��f��2��6�S�D&�����q�>�BV^�|�d����ΐN�z �,���dE�48�C����Tf�*�����	Hd]ȔM�+������W��W|��gΠ����<�(x��X'!��cL����Ď��UI�L s�*���wa�$�_:�Jc�0�Ad�j�46�=� Y�'O������Jك��֞�5��1��K�[.�Ɋ�0�0��f!nh�^�
~��]yh(���%Π∗V�P��1�Ǒ5��!�Ov��]���Ȏb��R��嵴_�˄��4��|E�<G^�+V����8-V���Ѱ�\�c�zhn��?^���c�_�.�,]ѰY�
b쏪fZ��B�N�:;�Q�p�l�".�1�G	6�>�T���5@�8��KF�'�v�a
(?�PfʨPO���X�s�I��<u��u��K�+H�M�NJ��s��,J������U�u�7��	b������!m�M�Y&<�P/x2���;o@�v_Z�*5j̑9��\�e���E+Ҭ(-��M;�Ň4@ߋ���9�~4'��&!�;��H|���sP2P��,y�R��H��)<��a�Uͅ|��B:4d���1��b����'V��d���Š�N>@A�X4��E0P�3`��`׿�S�N�sz�Hv݄~��Ë��(~U���g��;������5xF��f��V�l�"A��є���-��Q$9[�f1�|x��p�׈t�"���NV�Ew���+����Y*��l��̾_�c޻O3�]�vg��V_Ly+OS8��)�t(�$�K!ޕ��.n�$��ŷ�zV%��[T>e�q��*�B�v������MF�G��,��؞k���]Ld=)OM�|��=M����p����������;Dn��q4"`O�� �1��g�㮥t�ċ�<ȮW�̽�p��Xܧ�(p�xjE7+��t]M&o5��~��"�>R0�m'J撵�2�e���Xz��GC� ʸBo�2����L���?v����i���V�a�&�]Vh"�+�AT�@?T�F;�$w%��������h�h�ϰ���L�ͬ`�=kB*"66NvD�Q3Y6��������Q�9�µ����-s
vw/�^?�`l_��I�����|����t��T�ʉ5U�E���D �C!I�F'߀���w���e��ZSU5$G�d3�@�4��@=���(p)�G�ܥ$Dn�
��&������,�l;�y]GsR��q�f�V%0���8�W�v#V�K@�m��^�{	�J���'s([#V�)�������O0Z��&�G�I��îԪ��i������]&�I^!^ޓ*�C�/ֺg�1����3X���}����/��+>��4�B��h�r� � .R]J5fJl>�������ِ2�Ģy�����S����Z_hD�p�uP�ag��֖�k����S��)r1�	}��گ�q��/���g�P9�#1Y!�a9���޼Y�k�s~F�MP�_��/��#�+/IL
�2-������lU���B��-7�pZ�s�t����9��<餟��#ה�l�vG���~m����%��Nn'`��Ua�Ԏ�i���n1'��o���v)����4:�ݣAE�% �"�Pv��x��>j���A�jE/h���1�菖��K#$��UEh����:}�禒^d������o��~��4�:���vɳQ?}�iYW�m�aj$�Xy^�Yp:����XG%;��pca�I�2��O���'�\���DϪ�gx��ٷX�S��U�{�r;�jĀ8�[L��7�nlp�3R�3�p�V-�E��^h�Ve'����gF�!��t�K�6,	�����B1���������0�HP��"nf�3���hu����u��!M���)jT0�y�z��vd
��8݆��{QsS7����<s�fJ,=s�a�Ғ.SUi���wݷ���leOu��8S� ����p�M�e=���_�B�N�I�����=
������GN�a�=k(�����%���� 	�����\�E����Zl�`�ȁDV��3>�W��/����4謾�7��I��N���4u��:�Ekm}I5$>pI�_�m�L�E�8AMC(�"|��nkf�"D�����dy���L�mH|wV�� �тr� � %�_؂��v6+�[7�([��u��IsN�l��oQ3�cV}߸E9ӏ�vxop�˸ȥET����i�6�΂$�S�ض#=�۱�E	��w�Nsߺ��J]n�>@r����O@0�	!m�5)�h%�8�����3.�TB�W-r	3�)Q7�`Q�v"�� �`݁:'��6�s	�C��~i~7�!���T��DH�������Z�]��:F��w��E2�Vm��ũ6�
�a���Q�x/��ࣔj\c���+B]V��B�T�������[�<�Т�O)#.B9=w�0�3`�O
,�	�+saj�s���[�UB���z��%�y3O#���b��M?�l[��O)����ᧅZ�h��A5j�� ���y����A�(�x�[�'���d�*�~��.��>�+2̥���4N8+ka��ka�0�UD��T#�����/Z������*�=v��GYX�#$	m��pg���l8q?Jj�r�\�Ŭ
L�X����bZ�8����A��[����;���3�S����I��4	g�#$=��4���:N�c���l�WX�hc��;-�	'C���*�u|��h�/�;��F�xE��WHT�V�!z�|^OY�&m_ѵ0���/Ϡ�J�x\^�8h/D�[��:� #��V?f�|+�Q��G�w)t)g�)=��?�Z6H�R��_�2�{���=�L����&g�0 ha�fr�(x����Ek��d��_T'}���u���7��g���IB��g��',]�8�{��e	CڕĽ#ǒ��599(�ܻ����]��_CȻ'���%��F�ee����p�-�ı��]Gw�
|��t����j|���8���BY��[�+��^����)�Z��l�169X�?�]8_@���������"ˀ���]���[�]{�h�]J���3��
������m;$�}\2��|R�6dnIob�{��l�� (���OBD�J�|�Q@�:�\��H:��ob0��5{��-��C�5�eBQ���r��SSJ��<ڍ���I"�C���, %X��8۵H`AP����y(���C!��{�
p�/��d*=�4�|�a@����:��qy��ط�� ��ҎN�te��A�� �
��PUyƦ�pC,?����
�E2�J��`2�����f�'>�R�叉������v@9���>�!ID�:+JX���'�:J�@���"�6k
l\���a�.�O����������AT�~��cӧ��=o�`j��3�w-42O
L�j�.?o{��O��u�]�r����j_�n���1���)c9���k��ྗ�e���#�3V���U�6��=!��t����ړ�GT�;��+B���c[���� v� y��h1~f�z���2��2�[��%����=�1�v���BA�̵o�al��F�t�<��@,�I�5;m���N�g`��c�Sn���=óc�`P��-a'��z��Hx�p��pm��0�J2�j0:�)��H���ə
�y���07�6
��0�Ӿ�d�<��kB�{��Q�'���{���A���$۞����9e`Nu^Dp�W�#�%BOU��S�p�}C��j�K�M64�����M��ZC�ܨY��9�D�����}� g1`{u��D�A!�,�kh(�d���D��1�oB����Y*��gֽ������/�D<�-�N�=�t���)�穳�K�U��ˍ"U-5țoh*K�����r��
�WhO4�O���ϷX?��WJB>(�\HF]?�X�� �ѩ�v��ʥ��}gt<8Q+���-Σ���ߏH#v�[�Hф\�,�eK��d���x�M�*ѷ>-�I�>50�y�IQ� `j�)���*` #b��V�Q������'��ԫ��� 毳u)N����q�<x=lp�E�mGi2Ú{�ꮥ�	�σ8  �xap�T�1O��t�v�֖�뛜]� ,c5������ƫ�x��?)��q��L���E����ފ����O�S`Ìe��:��c�&�"�N�#�΂˰�t�+�]���)gO���z�ڠcP��Ku��%ă�wLY���G����_�I�`�2��v_-W�U�4�����o�f�6U��9�2�޾�se���b�##��z���#	!&��Gqy�͑,��a�Яf)#+�%+oO���O [�D�U9��n�Rj{A�Љ����Rp�c���^�����.�)�V�B�/�F��,��+7���ur�;�jn���#S�o]���0���[v����u�3i�|�;ma��(rS�tfL�cI�;b�>���˯��Bz� ���e�v&M尿��#�bHCE�ʖ�a��hI�֪����m ��x�>� ��������;�/8�!t�K;I֖��ub�z��Ǆ{�2�����K��g�))�BZ����l��
������$
a&n\���T�sL�Q4eζ���ڃ���~����Ed�W�.s��UR+��X��������y��@��5��<
ƛ�G��'��,���%q�@�s�Ħ����*�yiT��1v����&-��*c���E@�b!�W�F\���0�#3�{�k_�ۥ����x4H��G�4�)M���oL����ɵ2,oǰyyJ�Fy҉6/��6Q+��L
mKX'�ޭ-�g������c���iƔgu�ɏ�y�[q-��_3:��9k���o�K|<���0�~3�a��1���	��OC�n���8��``��P���rQA?�s���U�"[ㅊs�̞�>�{*�Z5 G��;[�(إet���9CY4TU(Ҿ9w���J����;��$��:�p���-�",:a������Y�ݗS�4M_�]�EW�1N��t��Ъ�+ݴ�� dN>~)L0hmJ�n�%m�����ՏT��}���*ڍ�����m|��kЊ[�ge�w�pݍh5�����.MvZz�u'���5��U�P+5���.��_s��#W[��,%�Y˥��U9�K�!P���,T����>ᔛ3��a��5zөԪ�$��W�#$���V �pf���@E�p�Q��JI��{]R_$�j���Q�I$�S�oc�{�͔8�
)�E@0�7vފs5\y~�x�A�Q?�:�k�ۢfO�rF�w��%� -��iUY�T7��n�b}��O���,� _���#�{� g�f��9��UBB}���,��}�eg����a .�1�ph�������a�I��늛��"��[�jt��Ũ���?Gyr
���.2NM�j�S
�&8����sm���ҞMY�@(R�_�a��qޮF5B,�礛�*�rg�W|N�>�0�^6d����aN���~�RXW���Jj��w�����˕���qq��ˋC��Kq��h�m�:t�#O��B��o�°��A/=�T�5��
�X�����K�iL�qS)�'���o�� ��9�xO��%mJ?xg*��9B����F�_��1�j��W�b��Da6 �ϛ��֬EV�� �ULU�6�s���3�x�fE�l1pp�c�,��K��[�~;��*?�\�eZ�wp�f!���������$ZU�O�H��sܬ`�ds�+��PVz6K3�D88�Q���������)cZ8�_�	,�`��by�k#��ǚfQ>8m.�*���aL��-k��/�&:C���E,�EB_�#�W�S�x���6��Z��`KE�\�o����Ԣ<�>��|z�Z'���Ӗ� ����Wڥ����ݻ��^���3|ǳ��9��.�̞\մ.�n�Z+�,��$,+��~��LG�B�2��<�#o͓>�~�qۤ:ʀ(�9�%�Ԥ��'4��G�R��x�mk��%Ay�?�?)>�dSs�� M0����U���EJ5m�MF�0%_��*�j(�¶G��@�2ʽP�*���,���/*��G}8q#����|ѝe{ %,�[�x��2\MR�� =g���)��P���݌�ES)���a�aY�@�=�04�W��إ^�A�& �_K�4]��L��.,��~���L+�j��<��Z��.���G��A��kǍl�?����
Ċ �b���
���f�5�jx(`�tO�z=�L���ku.�N15��_���,g��Y�[���ݹ�|�F��i�˨�9]<wT�e���F���}�&��ײ2�����b�b�w[+��]F�ތ�Ԏ������H����^�kV�xӞ���P��70\��	?C�Z��;ܞ�E����%ǛQ ��U�o0�[��7;��;�F�T�.,�70�N��n(6���Ƹ0���cыݫ�ɜRC�bm�u}0J�f
�.�nn�����t1�7&ur3��� ��ˬ���@�ya"r����2��PN��5���#c����N�β۲Dw��X`���f���F�#Xf�>��W['�� ;�iK�W��W�