library ieee;
use ieee.std_logic_1164.all;

--------------------------------------------------
-- Controller for testing purposes
-- Add components as they are made, so we can test the complete system
--------------------------------------------------


entity test_controller is
port(	
    clk: in std_logic;
	reset: in std_logic 
  
);
end test_controller;  

architecture arc_controller of test_controller is

    -- Component declaration


    -- Signal decleration


    begin
    
    
end arc_controller;