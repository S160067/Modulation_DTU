��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����0� ����遼�6������"���#�{A���'j�Qj} �}xT	g��F����a��f��洜K%g==�Z���L1������bG����XB�k6T��w+F��3r1#�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv ��i��X��s�-�Q?F�`Y�������� I֏�׋������H[��9����ۍ: ؕ��6ж���Q��" ��y&���Y	6_���.���M�ݟ����k����
۷j	���`a�s�Yot1H���\�GF��u�Hs���J. �J0b�$�e�SO4��ǢSIKiԒ$T��`�Ƈ*����C\�>�)'���@}�u/|�������"���p���n%�m�q_ ����=u)b)noпd[�'<B���U�N��p۫�W�h���+��P�=�kuH%Ҏ[(t)8*$��[M�,���-�n"�����;=��&�j���Ҵ������_
�@<��t���hP�7
����'NֱB��!���+�������@[_r���PPW_�B��U�VL�E�u7����3_/;I�.] <�R�d���h�Ȃ-۱	yvUШ��p��I�V㈧]2X� �Ȕ#(wkrjr����aA��3	�O)�H��|e$�$u���!&h�������(��{H0I��,�n�Y�G=�����ȴ��E��a�V�h�p:�рi�$:�;�I(��Ѐr�r���n��KOw�ӴL�~��t��E�A��(�i����~VUQS���;뮇��@�Zh@A�W�B��aˆ朽�6��x'P8�8��xVn��]@6[ymtG�g�/��%��B�*)(OV�4�s���	]k�{z�O�k����d�3�=��#L�-���3��9ƹbE��f�rgb�6�$��9�.��S�%�����#��l���Ԥ_�,sI	����^�	+�����/�r=��W��[�e���Aj0đQ�(k��P�P����X��}�������+�j��-���&UU��:�%ig��>a,�%��C\G�22�+m��`���}��,��ۍ�J�c�̀���֛���~�����$�c�IQ4�>����׺_�x��y�K��e�)&��"�g�}e�Ɨ����:�#�vq��m٦ڪ��0\ϲ{�xP�7P�}F��L@��JMq��X���_^u!�'?ӡl���{:�~�7��4��4�����hz-�Rɓ?��c�
Ŋ��[����/�b�;�q0D�t\��HU�ă��E�F�@��SMn�Ç���o��	��D	��sOs�"K�{p��Qn/�L��(%2U��y��=�Q��+�GG�	b��.Rf��^�:4a�y��P2E�p�h�����P���t�ѝ8J�	��yE�a_tYyvO~��4�A##�����+I<���ʁKL�HM�ESܡ��e�-��7�DbmH�����LՐ��9�� @� �Ӕ�s4X�l�>���i�|v����[M�K�`�N4m��B�1�(H5�x'��w��$:>j[�o�l�T�{�4l�/��G�|8�u��%?u��=%����mE^4s��M��սk�2�&�>��U��pc��@�D4�s6ܖ��@���E��Y���L?}^��i�#��23;���-���p����˴��=S���
)����fC�2LD�c�S8	����~�����{0Z�uQ���-�#�*Wd��$� %�X��=_6���B�溟H̩)e��u�H�+T��+])!P�x��"��������+�#��ûJL����1�N�	Q"C��W��i�1�!����|��o9�:*��{΁;�8Di���/�����'����Qv&Dl�+k��
Y&��P��^�]_�StgZe���ԏid!��"� (@��/�>�J��D�-w�!V��H�a��r'�/n?���#t`���x�{�o�����Y@�J6��]���c'�NB{��}�~���k��iDQہy(���� ���ü|����Ki�7�b��m�
�p�͌g�(5M˵ia���x�Q�P��M���A�a���^�\\ �7�twt���hC�j�=��w�*�2�K'�F��R��Hu�%/���њK��;����!��U�k��	�05�g�^ȁ��#�U�2�� ^�9�9{�i~��E<t�v���R>��-I�}�rf%n�Cٵ�2Y`[��1Φ9�1�3આ9l�)����ҁ8&��J����E"��9����Wn�P��C� �~����2�t"�p���3���xv�k`��^j���;�WT�.�l�-�z͈F�MY���'�a��`p'�ԍss����~g��me�H�`QU��푃x��פ��ģ������݈��K��Dh8?X��97��Jͥ"g[�bg��H�������r)"ޢK��.����RJQ����An����7�K����:B7�2o�UjAd"���il��R���3���0}� ?���Kۼj�G�o*�#�k��;��//� ��k�eV@�A�?��Sv I���[�n%�s��17gak�ǔJ�K��xV[47��y�A?�zk���K:�eS��S�yA�ۜ���1�r`�3P �a��x�[DMȱ��n�����t,�e�������a5�M���5��(�f6�j��A��&?�x��ޔ��9n�}���^Ս�n��%��r���[��M��f>�E��I{���j���j�3˭/��5�_�찛�o�Cj�f���^I�'
�5u	��U�s��$�(����,�[������ݰX�XE�V���w+Z�v��6�'8|�k�5�� , ��J��]P��=9�TkL��	8�ڿ"7$�p���o3T"�&�e���idW��o,��@}��.R!��g�N�au�G���Yn���f���dW�`8[?�W��퓏d%G�1���w��ZY#���T�Oh��Ņ�AK^��P����
����8��]�>�Y�	f��w!o��L���]V|�xW/<�"؉��
����
���饮f�쫈WKe.���}�Ֆ06�������[��G��<s/n�䖉�&19�8�A����f��2 (V���+��q*��u�4Q�uG���Wߘ��ߠ�J�bޯ�ڔ}��籥�M���"\��qGuK�D̡e�){��菉���TZ��hF-E����ZB4Ɩ��PU�{�+f�������O���w��	���=�|hL���<Xkٍ�����z^���`�<���3v��L_�����SD=���)�W��t	�5p��B�)k��cIq�i�%Py0i�=�"�`!���ʠgG�7,O����*o"6ÙY��Ǜ�fʽ3
{T�%��r �+�>��cH�`�~�|*W:X ��5�����e5{W��l�v��W}�w`���� ��=,A���{�����]�"����	+�vSW�&��
�UN��C��G��,+��x=Ca�S��F�g�7�1-D#0�eB��ajN��/�rv>2��ɏ����L�
���C_?~�	�-�W5��	�.���-x��]&�Y��}����K�>�?���Und�'�+�W/a��K�D�hSI����oH'U%�!����w��I�J\ڠ�	�Eg�3I���/e7�4�(��Hi3o��S�!?�.eS�|ssl~��;�h�fIN�n�Z����Ǩ�)�Xd�H[�@24�����4P{+��as��93�юHD}DJ�6�V�����c�C ���Z]��?�qYj`nz������u��v#�ta��у\�1�Ӏ7���f� 湑D��t��p؅�t���`�����Wݘk����Ac�%�]ZW���D�s?Ɓ�����so6q�6��&�y��b �s��Nu���Z��I̔��i�d�t�6ƿ���ˉ�w�1BNAWL��e8y�qiHB\���4�l�xw�){��g=vS/���3iH�������߈�A�Y�����'f�����>mm���<+s\#s�EOާ����r����p��-ج��KI;}��U|�����Me�Dboן$�>��y��qr������<A1�2�ʦ{p��Y�i���I㕎<:?��}��8:%G������b�a�ԾD�MbKuʓ��u�~
87��MŦ�k�\�e��BP�*��h7I��n�%�����L3Ɨ�.��Y���M2�����#�ߌ/`[�)�h��^{R�C"�bQ��ډ�Su���}�8x��Su;��D'����Q*[?6kH
�Rz��)��v@�T��d<�*�Ա�D��U�|��$�:I��6����l�q2����T.��	����[m,�o�G�>V#��rY����Ya�~yƴc�@)<i�D�A��ڷ� ���
�`R��I�C	��B�����fذc@��V@(ih?_���g7E�T��;^JCPp��~���(!�P�����(��R�th����)��^��,8��H��ϔv���ِha$�飲����m�1�!�4��	@��������%y�\K�|5p����Qkܕw����7A���v-G8�R��Z\��SYp\���b�}JE&���;�u��t՝QI�6��k��ܮ�%ջ
v��2��}TSt{�������:�r����J�ţR�r���$XZ��x>j��AC��\����ԽQF���0�� _��Me@����-Tk�bjo��B�����mʥ�7љ70����P}U��2�;�?GZ$��u��q*8�۝���5�+��l�狛f�=Nڎ�5ܖ�� �`%�`��I8�=+�n���(�B�{x�Kk 4f�؉�A�e��n�RP ���L����i�UjQ�i.�X�E��<Q��@��ie����b`ľ�Y��щ�ӜQy�F/)��I
V��,�שm%��f�<O��PܺS��Qt����YsUAS ��&�i�o�(��lC}��<��)=LP�<��l9�C���1�HA�C�?+.���SE�������)=����ѫ��M����cܜ��e�渐���\�c(�ع�z]ϫ�H�d���M	c�;�V�o�9A\�䤂Rt�Ízok��
�S�b�|M���`�{s���4���9��q������V����uT8{T*kxՔc:=��\�πS�)pa"ј)�}�K�r���{~g�������*�KZM�cD	w9+�G��q
d{m��3��0V�<f��j�����>4h�PA���ݼ�`�4<��gZ��u�b�pyI�0�$��iOZ�������S���b$��u'Kc�E�2�V��Qj���}���뇵͆��^�pݮ����~v��9v�Z��c�w`z_�w����#6���Կ�vG���Y|I��Hï���@��L��M��7���s��v����M�b7NE/�����έ��<�B<��H����cl~���7�,��� 
7	��{Ms)��A.	}�g�0&	P�������!���S��_���r� -�wr�*\"��n~��<��[��\����3�=KH@e�/�����1-��ξ�����39�ICX��=r�����a�P�4p�w4��d�gWƻ�e �ɽ�� :�G/�PY��O��V��`
_�H���JB��;2��(\\��u���ks�����A��;�W��@FV����3̌�P5�-��Q8PÖ��	��z�� �[����B;�(o��&Q�U1Rw�!�-%�e�wQ�+��#BvcZ�ן�Xy���+�4 L�T��=CsO�4������$�"�^<�RVx�)��y�����e&~�ۈ��0�kJ�� �B@0	�Xw"�i��O������
�'C�*9��p奥�I�%�>{z��!6tU��q���,��g	ᔖxe��X���ॏ}��G9s��`:e�6s�3C����*��	�Y�Lʢ���Vzޅ�2�^Q�,`]�lsb�� o�F�G��B2N�[�W~�^�{�LPU�fz����S��E^w�	�b�Ъ�)�خ�Hv,BlvK����QB�|�<��r�&r���+s��<!h�p�X��)�N8���H/M� �O0v`ؚ1U�Ʃ��
o��яho��KF&�%o$fه���mi.l���f��R#P
Q-���ײX��3�m�a@jF�;�%KJVo�/ވ�H�ot���"'��+�����g��︠ �i���`�y~��{�}���MQ���K-|��$q�e2q�:�HT�	��<��אκ%x�RG����F�n�ܪ"3��e��#Nb����Nw���-v��Ճ�km
Q�]��(����-f<뇭�WM��R����r��֨b���T�����}/�ŕV�dd�eͪ���N>.�ǳ�}?�*ҿG�,45��uy��j�Qh�ǚ���&`>i~��>�( cZc��U��Ce��ի�v�^�O�D>�q��g�#�E}�B�U�-�����aDJǶo�j$ #,�\��I�C�Ա���X(.�i.�+30��BXJ�?������O�A�r�@n��>2���]�W=�:f�D&�a�����>"�_pC?{X[�~gW��
��+�;$�7e����{��Tur0�M��X��*�AA����*��L{�S@��'�7������ŷ��M!�� �M�� h���i� P�}��*�y�'��0�Xp
����;ߪ��M�v�>:�.|oE��c�Q�)��Z�e�R}�� 
��`��D��(#A����VN�|��ir��@��x�!�$����!�8��Wh�-�1�eLc��q�H@z}A.�6��O�h��=�
���,���`WE���A�b�څ8΃���܎`��@��ꞵ� o�1RP�|8�f���7�?��HrM��'��΂��%\=��
(��#�,�a�p�d����*���`�T�N�1�(y���2�r��1t�Gg�����U�"�%B�Fe���W��e�1�R��Wg���6� e��M��M�.�D���!@z?T=ġO��J�x|k�ۜ��=��n6����U�����Oc�r�6���]�D6�+/1������a}��kЇ$���.)�(��閸/(��]��c�rX`9�e�����*��p<��^�%�H�Q�=� ��y�_�p�~jc+��4G���	��}�"�Ɩ�g
�S��#2��(6\T�f+$
�I�Щ7�:����@1��h6�f����iM[M�5Zgk��}���+Dn�q�",�lfmǺʇ&P�
�>���K��2;��s>�:r~d�`* �#�*p>!Nl{{�V����#�& B���7�L��3���h`�Hl�m��i��ȹ��䱨�|����Pw���B��_w���)��I��ɨzi�s�e��8�~1{7Bq��@rﲾ�o8��I�KQ�Z�Xp�&o�4���Rb5�ɏ�.�!$kԔ@⌃<NO�����6hR Gk%� ����fQGPG�6� ۂеWmd���\?6Q[ȜM}�)�	Sd8�&�܇�4� �{���2_�y���2՗�\F�]�e��dz���0����v1��+y��z'P��
Lo��ӷ����	u�v0xW��X�A��\���G�]�%��O�2�]��ʞ)���J��9+)zmp�1�4��	!��>��m�c�ڃ���#�9�� ����mP��R��|p�M�)� |�ՍZU��$�g� �/ad�@7c��6E�>�j����l*y�?��;����0h��u��|��t�X�l�	>9b]�[��ƪ�:Ũ�"|ү�X�6/
�-�aYJ��h��0����9�)h��?#���V/[%s+O��H�bw~�~�uNE ��_35F��т���(�� �2��O�Q�b�m�QcMC�O�TssGr�7�3SW�,v��L8��S�ģ*#VZ\�-J�[�t���}$V/��H��DɻW�=�`�%sc��c�F��\��Zۏg�~�Ggźx��C{-Ĺ�mq�۽�|���~�լ����ιHD,@�| �~�"�"B_�}�i�>Ћuw��R���{�:��H[ڷ��^{v��/�Z�q��y�L�����61cc�3&�Ȳ2k{���]0��2qe2���/�&�Z����l��Щv�~�����р%x�@����q@�{;��ߨ�g�r�7���5v�� P���>�B1jL��[�{U[01��=ר��J�5�[�&Ƚ&������������縷l�Y�{5�^�%����漖�8_��c�aMa��u8��Ơ��ת/��g���Ct���P�qg2�d����#���<��
��c�ݺ�tD���ܗ��bl�u��wĬ���-4�yV����St���o�:��Pد��1���ק��b���y<��4���.�i�D��Z~���{����<��SEQ��ʷ���J��ץȋ%��u!ӷ��?B��D�x�#꫏�e���1s[���l�	�^��%�JI�qE�♙uk��F(-w^'�����KE\�X����W:Z{%���O��}?/T*aD"�]y
��q�����QX:.P��pbY_Ol ��%���шM͊��o��p�RŹ�'�S��-&�Ux���t���(XK���{pN,>ڻ� SDq�F��td�߂$�N�7�����S^��p�dÔặ��Z�	ˢ�_(�E��s��m�O���?K�8O|Ij�Cw�h�`@v������$v��i��w".�z�`�������x���[]��䨉��V5@m��n�c֓�V?���#U^�����"���Фs�3�",��۩�؄����yI���,l��i#����%�q�H��6G�`Mek�����|��F!â�ر��әf�q�H�o&�W Uq�~~G�3���f�J�m�2hgA�\秭�����v���M��K��E_;���D�4}����A���
 �a.="g�2j^��Dog��f��n����3n�?$-��&&�*(\R�����|���m�R�urG��3ȉ�!�?p1����Aw��y�C���v���ʥ�C�?�Y���H��.�e��<ʪ�$��Ɛ����-��#�n��z�{�S�SUƩ�[��^WerͰ�F9���]���V�-�}7�x���e���n2��~ʵ���>:AI�\F�f���A%�Q�;�B�|[5)Z�tn������֑(��q���J3�Ѕee�Zm�[��� Ć���@Id��-�Ii\�՝x������(�T�mk�^-���(�#���0U[7�XZkcL$.�Y��F�u����!$��cw��̫C��{궗��6I/̵,cwr�-֊g��5��(���i�4����M4{�S��N���yJނ����}4��%f�*\	1x�FGN����E[�j�1��b}�W�=I��x���'e(B[�0ṡr�������4�+QY׫�z]D4��p�����u�+]'O�W�j���X�5�*e��Q{/����7�Ӈ�e�,@R�W��c�bg0���q与$���]H��zN��.�طy��$�#�6y���Ts��p�*l|���3�5i��J��-rz:t)���ז	�e�K��J����{�Ȭ~��D��ޜo1p�V�~�֞��H��K�v5��V�9 ��8������$6yPn(����V�u��̺ӯn�Ș�8W�Y����A��6�XC�uC���B�9B�̪!gHIz�s�J.�H�P|YGy
O�#�;[�N� �ݫW�x�:mB?���:����
$����N,�Lg0L6�:1�ףV�N��iG�y�B!X��)O�˝ը����S��ש�ZO3ؖ���P#�e��ی,	�i�s��0!K���9�h����s�&�U��I�A��)E�����v�-q��3�U���c2n��"̘�������CSYo�F�5��%�(Qp:8OE�����A�
R7�q�X}Z�?<��t7��\��J��<o�T+��[����8���3Û$�>ع��P�nO�cy���?Xh%�o��%�U�a���5b����>�M �t6m��E�0G�-<:���(U/&�{}"#E���M�vd �|��k���0��J�.xqw��$�;�vJ;��>6j7�Sw���/�*B
T�0V��*�S���e���4�DKdm� ���n��<��>o]pÈ���,R1t5M=�~ԓ�Sj�P2�`�N��c�Q/6��A׹_<,ė�! 2��|��R�;�i�R�#�~p���2U�nv?�b?��PI���qZ0�(��!�MC�`@cvA�G�!�����[�1f*Tl�[	�#���7c����MR�6�|*��]DɭEA�.��������b[ch[�<$7���f�j'ɲf��B\��FN�>�$����F��^��h����S��ƶ�� �^� ���9!,�^��'q�Ӫ���q�
e6���^݋�y��p@��H�^��a�#��@��$E��SOZ��ʁ9ɉ��OxW5 XTQ2K��\sRN���~�8�cGߟ�����7Z�qFޛ���9�T_b,3J�~����j��ʂ翹N:;'#2]�@�`-�^����<|�W�uIT	��A� �]�1�r����!�R2�`G�_?�����ǵ>n'�Wv�.��K�T���-|����w� ���� ��n%�T��L��,���84��;��a�+�]���*�a'��C\sUj#{8�Yt�k:�B��bUn�o���1ڻ�4�5�wP=puǞd���c���^�׹�g^	j1E�e��q�S\��^�9��I{1�P�%@������S6�©xj�e��f�ꑪL�a$&�l�o�%���{�G���1
߬&爋�CM�q,n@3�
>�������fe�{T�\&B����ňM=�����FA��;��{9\Z/3�Pr!�I9�6zН�/�M~�����	�a��P����99���S H1�R��m�)�^�^n�#��qnlD�a8���QQN����N��0���Pm?b�e�6����]	�'��hI�����WÈ���G3o/fV�,�nE?
� A/�N�	.[�@���\bG%�V����rCk�Z��x���)'6Jz)���Ǚ��^�t�[=p�5��@>Z�?a�ĵ@T�{Zkw}����ah�kX!�W��QJ)t�\�N�B$�it����G�ޯ�K�i�M �����f��Q�-iՠ�c^��ի��-����Ɖ�c�^Y�5��bOgyOYfO�aw�&0<�J5������>��MY�[�N1���-�h|�Q>.�����	���m.XL|�	5,|\-�c�;&�ß�e����t��P
/,���p�<V�1�O~	ҙ*�=�����!��M���T!����*s|L� wl��_�G��FH�{�Ms~V������(6�I_!��@�M����SNِn�Ĥ�šlj/�7@�ӂ4�_��ބ�E�m4U��E��ߜ����5>����(�쿂̀_��N�9c�R}�����"jY�l�s���x�Ϧ��
X �|�y�Ĭ��b�R�j�x�������yN^X�{�E�1����!P	s�8�#��Ew;�i�g*��"-��l@��q�̘��Ux��2�Zxʃ���R�Mò���p>�'����A����<�ޞ��W�yJ0��	���~�Zy�i��8	�1�%�@�Vy<�Y �V>C7�S���)����n&���ڎ��)��wb�圝��F�9�k�M(�c���W��]�����W���N��B&�P.�	�c<j�cS��[�5`r��aBeA*�TGB.��K�ٟ�q� ���RN���xk}������Vb�޾i���q�?���!��V
]��M�6�Ny��)@�,9��oe�&#]b��j����=<�!GH�V��확�I���F���"�8șӲ�8�P	W?�Q���c�%31f���'��"�Y�ɸ1l�|�R��n��"t�O��Vg4TԠ�}�	+1�#��R��fs��>@e��f��4�n�W ���+H]�>/5�&2X7�����Q�l��Z;�̪e�RَnS��.��;��!vB�a�7��GL�Š��|����9ڕ/�b

��~Ċ�Y�'	tj�.�S���ѵ���:!�.wQ5+����Ն��-=!�M'�!��dSj"|�Z+*HǼ�2J�@���iu��x݉h�����x��h�/sO��5ۜ:��J���c#��8�ukÜY[
�D;�N�)�V�8�Q9����G6♒�P�YO]`z��!��@���Ξ���j<���rE����l����E/��>�~ً��U�~p6�K��#��,&D"���3�˰B�ۜ��K����n^�Aj)9��mP���s�yUk�{ %n-eL�l����Il9�inj�JL�R���AX%�7���{���\�e��&P�"�	D��	��ON[L�+~���	�Z��@��nԶ��Ru`<z~<�i_ND��`���4]:����m=����ɨ��ٿ3
 �R76=f����%Q�M��R�+�3"am��F�Je�D��o����)�M}��t4M��O^���/���Z(��o�u�玵�f�r��.�J�P�1i�Dk<g�a�n�� gyzI��}ke�4�F�|��Y���[��@.�y|�����Q�)rV3��!�BO<��F.�I�:g�sjxƖb�u�6����cn&����(}0��7`�SQ
��G���04W��|T�u�f�R )����#~��8$�˚G�UW�RI�'���D4�Al�:�Ts��'��6��rg4lV������(�$���h��Ô`Q]@�(x�aE��YSh�v?L������w��8�֯��<$��M<����X����{W�j���m�Fb)�k�)?iY��`�]@13L���ti�J.�2��B�c:ч�"���a���6�_h��?FhXZ)�e0h�;C>��ݡxoPUf��T݌P��PgY��pOk!��6��kX�\cet�`���2iRg9>���Y�����_T��%�H#Q�����5:����շ*h��K��6�>�Y�'��V�sƒ)�
�8���7���$c�(0��SDA��
�k�+ �0t�u���\��~&���-ˈ����j�1h�@��}��q�g�:���H�ٱ]2/T����Hp_��YT2�ʇԤ�����%	ꆗ��Ć��J ��w(��e�-����|�|���>����	�pQ�5�� ZK'���'��>%��v1ٻ�:F��͌Q@��-x�6�je���>�u�_^�-0l¼.?z`������Q�D�x�E���e��k��~C{����E슻ہ���;M�B	����*�S�?����}����V!���b���K�� �xaS���j��b0"`���e�|����*e]�P���e�c2� ��J�c��O�g��	��a��� !D;����Gs.��U���_٩$��fЫH_��7�:��X�� �3�<��8�#�J0;י3W�C�l��f�{��VoBH����Fԏ��5s�g$��PH|}z��ITY{��m������^a���9a�������+�cn�/6���gY-XqD��1�&`���/��,�\�e8���xj�^*&;"���<4�F�i|�Kǧ�?�|��m��j�gE2���7��F߇P�"K��qܜ</)��/Tq/��̍���7k+R�D:��Y��`H^u��J�7ݪJ��������ַw���(�Mҿ����Z�Ud� ��~~��� N�7�CNV���q�aM�^����j\;+_V���~�-t��dMIͲ^<��܈�M���t�1'�3�P��x��g+v���� �SN��T��f0RP���,��2���A^F��y�ɺY)1!�Z^x2�B㞹��0�t�zY����6䠴?��I���/]�o���g�3 ����r.{`ED)%�"mU�{��a���qH����"���4s����)\.��~�u�"u���ۆ�|r!t-�������X Tn�#����>x}GҒ�૙����9�������s@n������B�*�y
��'�N�`-�t�W���_��#��t�\0u7�P�IF��L�I���B�=rC	���n�W�m�@���8'��r�~ �o� �������[��C;V��N�޲n�v��2����qz�2�$*�\���t6P���s�~
԰�*���K� *S��f:�KG�X� ��$�w0�M�O�O^�4�_�;�6M�])uΙ'��g�C���/'����e�N�����C[�b0N"��P�9���烍�!�9���m�r�j	l%II���	m�S}z��B5}A�q_�'f(�˾�d�.0��
�|l�$rKS<��X�t%&��ܮ}Z�8����5��U`��v��b#���If�0���6h���5�Ng�Ƅb�̒�0$�@��c�|Q&ѡ�ˆU�PH<�^1-r�J��x���������9�I�����W/A_;������yC.:N�����,ź��d��/�����Q{���hy4i|���x\Uz��w�m}�`����<�W<�v��="��f�eb��{O��)����sF�S�@(>�=X��Bt�_�xS'�k��=��s�%�}�W�r��J$�~��|�;U5�e�u9揆��>E�/�唣�!~����m�gVi�ԣ<+(�y���g�����J)6�e�����W$i� ��BmB :��i:ҸCNv��x�W|-Աw1k��^5'��è�m�h<���IX�o��>Lq�{)��7�J4����&�M�p���T����n�ʋ�aPB��r�
�:mH��"���4�`04BH��hρ�7���
jd��I�ƺy3���}W�I�>�p_ߒ9��Ħ��`�X�+�c�(�A�e�5|�;��#l�8oݷL�kr���� ���ֶ -Z�Ú�M�d�޹A��V����W����*�s<x�/1��
�
���<*f(#�Qz�#���s�^dϿ��f6%��*���o�К�K/�?-o�W��(�xt"�<ڪy���FHV~�Z���߅�%5Z�q���ԃ_�G}��{?5HLu�����[�����~�q��b�t��X��!��c2ID$�Y �ȳ�c�`2�[����r 9�>��]_� �c�-�I��X��B��DY����Q��3dA���*���C��?�����d(�˲{{y��ڊv���u$�{ʧ�mdֈ�*8?�q��!��4�	"��� ��$(=����|H��H�N���ȕG��A�1��&�f}r���.�#��g�"DU�8����x�ˠ�V�H�^�af�1��Ԛ��~k��[|�M=6�����mW}��%9m�ZN_�>M�Ғ��	fP2�����Iő�T�R�11mS�����ƞS�b�ῃEH}�7tWq�����-�d�:�#-��dܑ]E����J�߯3pD��#�)�A�rᏺ�t�c{�`��6�Xs��W��u���&ri�:��%���X�ޥ�ۦq���"h����[�����v0��'6��g��Qr�z����q!�$�~��\Ҵr��kX��> 3�.Y�&�mO�ײ�U�M���}�Zm;ڗY[�hƨ����-��^uW����&�۶f�4�1�?{�}5sI�������s�6�%8�>i?�P��ub�t���ӻ7��&���v���W�xǦ�g�02M�i1k���)��/{��"��)�@Ipٔ�����kA����ylg�㉻k���-�U |�KZ]9g?2�̗�~z���0�l��P9�������T����q��j-}0n����jF"j�Huҙ!�����z��q�:na�������=�-��:����ɠL[�/����TR4���j�
8	P2@����4(��|LgP�j��t�����1!������b�Y�|��vͿA��P�ˢ.H�/��jA�d$R�� ��W'd-����VG�m��,.��>�{G����r[F�r�*u��{i�I��+dg,�]ӧ�'�n����� Sg�����-�Ũwe�QoYA����]D�t&�2���D�R~���+
�f�J�OҀf�w��lI�1�
�ȓ�H�{��d��/xݟ���%��r"���0�]3.�2/�pm�x'J`�U.�wÂ����t�C_5崀��u 0��=#��{�(w���C���B�L�騫�Qx���za���#�����f�3�[�Pȭ�uǳ�ČܯPZ�-�a��C���c��W�J�k� .�[��+�2p��dw|�|?ctM�~�t=M�R��s ,��#�)�8��+}$�����1-�U�M�Q��tJ[�;��Q�xc(��5��dȤ��<�{�� ���Ơ����#�l&d�]C�OL�R��_�D'8�:Hp�㨺t*���<�.��C,|�����h���U��T� )������G�:i2��M&y�b���������	�8y��נ�K����o�lb�:c��G����4Ĳ8��H�.4N�������\�S�5��"�g��}z�;S�>�_��B((�7�G�$�|�������9ݦ��>ss�r�d����Xk����V�����N�mJ�<�!�C�(���� $�����$އj���A��e�<4NXI�o����#I�z�a���p2�<2]&�8���ҞL@�~,�{.V�9�us���ƃ�YH�6Ê�'�6���?�*�L��?��	�߯�r�%��rt�T��4�Ά{~�`���kR�l�L̹�1�u�]���V���Ŭ�����q�zs���E���^�TB�p���u����q����[B��k�"^����n��;PV��'"��K)���T@��g�j�����l���t6D�`����L�&.�O
ڦ����].�U��l ��?1;4J�ǩ�8W�hԵ�2g�h�)Z�~�����,���� ������i*�)��x3��^�TLN��ii�x��DD��*d0%{e�@��vk��p��?�Z�Ϋ#�.ٱ�?�;�b��������}�L[����n��v=��䊴�J�Uq&;��]u*%W퇒�tG��i���ͅ��ELTF���G�t~���ǋϢ�;׷��H�P2���ݞ'�^���{�yc�u��#��ʂ#��s�FeEl���3�U�x����El~��aiz�wFK�MMt�]޴\�t���������#a�����.i�ƸT(N�}B0l �/&ʸ�v���{����E���kG�lK�W�}����ǥ�/Qf53JF�_�K\��$���'a<�:�KĚf���`�<+�N��߀�����b�_�ͺ
@+B��9�_�������M��l�/��Q�������}��"H�Bl��c��4�'X}+�o����!�z<�[4�D�뻭�c�E��e#K^��h�Yz<��f2���&'b�vS�������ά�[���{ݮ�?����v��<�C>���ʡ>� �.�w��u��H���F.�:������_"�6����J[�A>}'H�_����Q�G�L0���x�4�tx���G����#R��QI���NY/<��b�[��ɚ�fXƣ@�~�J�7��	�褖���馅H�����	��f�Jqb�d^� lH�Blu�&P�>Q|6'��#���)����g�5a�ă&լlD�c>�U� ����� �������N#����V�#x�0�	���r�>�\�xA�lFz@+:v�A���U�aѮe���Z%`TQ��{�o�9Ӟ���<H�'τƭ%���Y�J�L���2�	�da9��z+�{쇄qa�q�|����3�#�DnC�8���Q��LAN3����kùDs��a�z����˔��N����,��(練��{)��V�ۓ�p����NT\T���#Cؼo˄���{��N�.���s|[*�)�h�
��?mw��_`jNۋ]鯟f�;�>34|T�p���,| k�3]!j�H�b`g"~ߓ��J�E��m ��v��~�W��=���a�Zw��U�&p��3Ȇ"��}g#?Am��i֦pcY���])8���DG^�巪���M��ad�o�f��&W��v���\ P��@ґ��x�^�e�rl{xi����V���{�7H}V��=TZ�������\�Ep���9�,��B�����~�i���$	�\;1Ϩ�+(�&�f0.���nT��ّ���-�}���e̖,Ӑ�B�V+�1��1�cjD-����!k�����@�ن>)�Պ��.i���U9��!,�卷G�ܴu����|�L�	�!�!zόx.RgKf�S��9D�������LTg:v��ʷ��,{�̣����g�\�>�:C���32L����P?��[ś��D��~%�o�4>��yՋ�N6A�A�nss}��M}�n�'��}>��X=��<�QJWr�]ޟxJ0�W��O�%A�w@�WU֯s��GE�����,�yI�I����L^C��LY����`S8G� �q=�|A��ߗ��R�ki�t�E�1RL��Jn��d{}�����᜚�D�\��yބƢ�R���>�L�e��]�|{�i�$��|Bٍ MK��?��-�f���]?4E�5�9Ve'����e<���Mi��ƕ�d{����@"��o�5T��f�����ޗ�9-�0qCވ�@ڭ�k3.~z/�k���)8��n\�vuy��'"����g�w�L�e�2$���*}.�|�Nt�^�r~�(ze���9Q�M�$�$A��E4�=�׬�ʹ��'%�^��ľ���b�V>��� �ne���X1�w6�/pcXJ������g`$�Q�U�(��Ԏ��9ӷH��֒@��t�X�S]�z��hR�6�����)�z"
C�W�E"�2��/���$g��͘<P&p ��[�2�Q�(˒�a��.���(��ϯ��\���m�U��]JH��Y:�o��vf@XbV�b��Ni�$d�Y.���
��1�M-Q,L�� ��=3�����YY����O�4騶<DZ�$L�g����{T(��W�._Q8�{3)��- Cn1?���q�Є���s�[
h��f�&5!�~�t�4�+�� i�h�i�tF��Wk����	#�i�B����M�bgW����Q	�G���Ϯ�x]��7Us �g!��=[g�&mq�Xa$�bBޟ�Q�������"Pr`OpO�8�"P0��$�y�y�'s�TS�g���GV�$�:�������++�ߒ�$�|����;ps���z��5y�v�[
Fԫ��Nm�9��j�P-�dl��T>2{;ޤ���Z� .����(����	P�ZϦ�����5��W���z�Ȱ�rOe��ؐ���W��C�cL6���yp�\�x���L�hN��^�~�BLt8��W�$d�q&_��"?�ֱU+͎n|﷔�V-:	)�s[K�σ��Ӛ�4�3C)�uw���Rr��`u�pe~��ٯuW�Ga�&˘]m����.�0qY�Q��W�/�Z�a����>����@��qQ�Ҷyd��"V��a���%�m͊��Y��\$���[��\hX���]F�@K���� 5�OJvi�?�AٞQu�|99��3Yߌ���ee#�"�s4�����=A�x�l��Q;
.��0qg"�S��z�����wI�^
t��pm�H�x◁E��J�M?u���ES�Men~8�_����^�;�������gs y�*yh�m ���;������+!b�:Ip6�%ř��="���,�F�|�t�q�P��\�U4���r��b�wiy^VBCt�<��@U���:���N&���5h[N�Zvܴ<�t�Xu-C�^�j�MW�ۅ� �[)�/ŀ��E�_c�E�-c.+�̻��=qv�� ��xrT�w��b1|����8gVE�"�4g��D�� ��l��:-�o�N� �����~9���SϢ������3ڃZK;K�E Pow{���m�丟c	^�P�G7�������$L�e6�O���O,S=Q!��]�t�z��-M��'����-6��=�8a=}л����?����m;��G����ͤ��&|j&X8��(��` �M͈���D����	�5��"�.�6\�{�S�����tU�����sk܅\�eZ��	���C��ype	��	�ng�jۜ�NX1�!h�M��^��D�9{o:@)����g�Q~��9- �כuw��E�:�/Q�hI��	�����G���Qu�U�gm[$f�2��[�p��ݘ��n�B��C3wroŤa�4fR��3o1cf/5R�O�d��#6�_}:*���������g�Gb�e=PN�t������᠀3g03RE�)��B���{�y���fo�SL��w������LF.a����J���=fEC��JZ
G���f�޸2�yxʤ�?���t���`cE���m�+$�Cd֜%��;�*�l�te��?�S�N����: T6'����s�\��6V���Q����g,4���Ⓤ�� �&)�O*���U� �I�ҫ)��S�����Z���*x����(0>��M����ВY���֘�ܹ���`��.��/�,{� �Ǩ���Ƚ|Ûj[y��S���/���8�s���������נ����e;��X���H_�;&�D��t��)������J���HUUM[�����p�ɥ�>��H~�GJ��\� @���(��ݑ1mV���7ě�%�.�&�G��"��!��+�h�Q�_,WԽ��ј������x1�n**�u�e���ښt|:,#LN�ǃ��k |���P�פ�)��pxՍ�4�L%�� �6��0�����4�-�������shj�\��v.F�e^0	�شAN�b@�]�8�i������g_i��7O�(�Nu��/w����ڹ��s-nj `�M
U�g̛g��֑_�i����k�D��-3}y����^g�"�\Og2�bY-��b�
@�X�9|-]%�d�����j��kw��C��-�V�P�7ݪId6AS��w
��=��Ǖ�A]sJ�M�2�<%�2K3O�\�{�B(c���U-7�f5�uіL�x9�QkŮ��+8l��`_�|�W�-O��D�����L�dWޔel��7�h�P�TIX�vS������E�ݯ�  4F �#���]xIkV�e�9v�΂��Gv9�w��2�s3X B0��r�\S��!����8&R���$B���v�A��W���G�d��n��ӝ��r���w ;?�C� !������{]���z��lTD.�)��f�ƻr��q�h9�%W�)P޽��_�bl)�P������ߦ����%�!�u0�_�����	��f�o�s�{ʘ�n�7ڼ0u`6a9��yg���P "`D �:"4��
i�{pg�Q��цN��[{�J��Kd��OAp]�a-M�f@��/��|�W������9��!�1\WG|S� �ƶ349>��u1��"��
����=<�u)��ӧm��qm�5$=�GD�(��b�(J{[;m3R����C�6!�+E&|�Zg~��
��ؘˬ�7�ҍg�dmc%ݔ�b{_{��aci`d�_��U�S�jQ��fq��[��R"�<9��!�j��5���P=��X�VZL+����r�*`��}���w]�Y�9L�|ձ00Q��$�5l�ʁb)�u��snq�e��3�9푂;Ρ.O��jl�L��
8��-�&\�]����=�g��=(����-M�0�c܋�A{�ʹ��AR���{��'쀊
*E�=r)+��k�O�}�.Zm�T��V��>P�Js�]2���
�u	����mK_�Ջ����~FeM:�<���e�!evP�+�6'�}����x���wA�Ǔ`;\�1�_����@]�
u�۩>��5�:]\-�#Pl`�8J�a���ӌ���)�W��2�,��Iu��1�vҘ<�ޢ�4�=Xr
�������
DE0,((ѻ��w+�pb~��&r=n{�m�
=D�1��uoP�z:��T���+��j!���r;&Q
"J���s�`�[���;_�-�q�����<Rb�t���O@k���Dpku���N�.���,(2���6�Z�(k��oT SkyƠ�shh��\�?!��)ҍd�/ZՐ��d,����嗕����˒Ur�ts�����}���p�vOS�h��C�l���t�4&L�L۔��}u8�a\�Y��e�'%6t��ƚ����׹)7!fԀ� ��<;ޡ�w��y����o�ξR��{ŝ��'y�7&D҆��1W�e�mR��+v}�><i$N�)I��sm}���S�����~Movs��6!�9=��5[W�2y�H�!f;��\�sL�,�����ԕ� F�*\`N�@�jM�Ӣ�̈ŧ