��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����>�S��fI#�l7x%���$or�#�6�y���N�i� �D��f(�:eǊ�` ��S���^�mBƱYjA���v�0��kh������#�v�(#W��ux��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�A���0>�kz��/ �_M��<-�[a�%�����'(�S��jS_�,��8��T�.B߫C|��N�(ݝ_l0fS!��mYԥQ��DF�S;���h/��9mϓo��ޗ��(����,n(酩���5�gJC����cKa���?]j/�a<��/^����G��P�T�ȟ����A�PJ��4���'��)Q�;��lc��'H����bm��9z\��䱻��Pp��;�$�@t��C`�s�7H�!,��b4�"m���!0���}Ɓi�<\�*I���,T� A*�u�
��~(C0�2����VN�Z7�|9d��21�57�(��v���b��T���1����э^���c���i�l	�A
����q)��vι�=,����S�ɲfI��E���j��Vw���]Ό.XXv�TY̘�%�D�Ą˫ŕ���^�")���p�����r������oup7R���3�ߦ�̧�Pd��1�_
�J%:��Lm�b���0r�,x����Q������@���.p����w:R'"5)�����@y�$?QVx)G��!{}ZQ��oȤ�ʳ䤬�Q���0�[Q�*�W�ɵ���������=�B]rR{bR|��6A�eb���̣���i�C	x�����i�'�D.��!u;�95�Q��ɯ�+��>V�E:?�2h4�������Et�mA�=�Ne{�)��c�up�
S����UӸ��G�CI�G_�S�$VZ�~{�b�/��C�KlEX�)���tY�Zz�I�`v�!t#Lf-!4}?D��g��> �r��	����|X��?�x�v�W+�^܍�6��?(���(�}{�ұx"a �}����7�ڮD�_��� `;�}#�I�(C&_~�T-B�;��=���ɜ�ţ�|��\-��(mef7��f��p��!�^�>��I�e/�+{透'�O$���ؾ
SOZ��1Ho�c�j?iZ�WJ�S�l�n&⋤n>c���X���礪s�B����5Hn?k��%������p���.oE&�t�q�K��/���� .�m�7(P�=��
m˴Vr>$>�Y��ޓ�9x
Ux�fJ`!��ͅ�Z�+�� I�1P>5�HW�զt�l��l���X5�l�F$�aoH���1�K��C��I;
0��|�{���_�gC����%��]�9�>�q��x^}f����0xtE��~���D�;�|zj��|�R�3�M�h��{U��"�}��=��73��b�5�~��2�JT�om���AT����|%\o��Xq�@��i�]�֍��J�=,BT��{�%h��¿I
m��lEz�F%�<�ȧ���H��*�zz'M�R0��YjN�e(?�?�
ⲽ��}5C��h�Vj�����d:�2��D���ȯW�&��n�*G������A�Rvj���P3�Jݬ�4s+$�~��i�N}��w��3 �:�L��ހ�BA�#ڗ+���]:g6�bS����b���O
�^�s-�C��r$Od�Ծ�&yd��K�_��"-u�JX����[���C��9��Z�
�%���]) >�G���B����H�_�j�[dd��1Gx�43��p���#�.�r/g��?,̔F���#núI�?�8t����4��u�l"���/4���*@?�2�~�L��v�p�S�`��kD��X��!���B^��P,����U�;�1�h[����/��L�§��0�ks�d���'�Wh|�"<,��)aEr���A,j�yM���3�8��b>;���Z�ީ���U��}�Q��g�mZ�gD'��F�ߏL�'D��+T!m(P�M�á��^�LxPo�	����) p(��D*@�k��YN�(+��n��Nd}��·��B~�}�3�k�f�ۯ���'��ۄ�l1���\�W�:������vVU��b 
��<�����v)�5e�Lp>w� ����X����h�d����5;N$���mL/juW,���j[����w"��`�L��|��Jn[lAR!|JKZЫ�B�?���w�
񱂀�+�;�o�-���Ƙ"�Ĺ]&����_$ݦ��W.qE.�h���P�;�d���g���<�Cx��z��k=_�ݒ0p �FO�����2�QL�"���� �tA�"��p�Y�GWZA��X��5lsX��H�ە�2=)?�mX��B�쇽�;�X��ڤe���Mu�+����h��:��J���z�`)�z'h�Pĺ4PαV���_b�c��9��6�zX�7�""�j�%=^py�����/urhB�� ��G��,����	�^�R!5���(?9�#���������$�a�*ʊq]h�;���%�胂P랙�ʿ$b!Re/������t����4n@��%Rs��B�jV�%��"/m���8'�Y~�
��@J��cQ�D�n��t�m��)��@��U�lX��3��Rnk?~����yy�6��w��ܝ.Z~%0z�����k �0���,���*���u�ؗv���JC���¦i�`r�~!�V�`��kb��g����5U�{#�I݇Vv��E�7�84<h��+m�������u4���6�{n�n����4��������狌r��x��(9�].��]�oJ�CL�KP4ʾY?Ri�"c�Պ��a��
�Z31��5+�Y+d_%Xzz%�q>����<�>�PZ�:��m@BO��z���1������ �L�W�����r�FC��я����S�Cp�Gǋ��̆�b��(�D7�|[����T�!�co��\_�;L	L���~"�c[��i��Yj�}�����r,Ҕ�����?HBS���G��i��=�5�}��3,M��w2�9��o��;�}���7o<�do�`��Wj���@��"'���BC=^Kh�2]����bX�Y��7(�����^/��FvW⸃Z��N�bo;Vb������Q�K�Ժ��o�̘����\`+/WL:�ԋEE�;��a�%A�KA��X�.�Qv���tI�z�����Tk�ڜM2����{1y��-N���z�,{�n���n���uD#�꣮���S�}L�}��h]Ot_(�KyĖ�]Υ�?g0_���x{O�����誀���NX�oQ�WztP|O6'?��Z��LtC�K�x5��	�̑R뱅d�9ӦF��rYxX�z,��R�,��-�N��lB;y�khRX)�僲��9/ٹ���g�k��X��
��Ye����n���Ur42CTcy���/����@�-*��V�i�����+ 2�`-��i�Cѫ��ys�
�^Y��� t�'��4%�6�wK�~ux�_�I�Y��6$>�)-w�QV����7���ǿ�9}���?x+x��m��M鋡�o"�`���y�_3����+1��Ǔ�^���'�\4���+�G��6�Jw��n�Euh��Q�v�V|���:.�9<���^XL`H���W�6c����wH0���U�Z���Q&N[n�%�ЧL}�"^;��G��L��E��G�����D¾�+i�(�����{ʷ����Vй7�M�~`����l�g�����4��
R�]g~��T��[Kr��~k���(1ng2��9/�+Ih�yHϏ| �؀Y΍��$%�#B>7"�"�v���PP����pQ3L2�9�p�����/�6�W�*�\��ߢ�Pv�7�99	:pa�T�1t%tmQ3�
�����I��sG� ����&�N��8���<�ǿ֬Y��&��Z �h��8���l����h%���}��-�x	��$8Q9Z�n���C$]�k1��Γ��@#v(�"%{=�[ 3��@�#��P�|/��7��B��a��Ѡ$J$�_J}$^��"A䴽ơ@SQϊe��	��j����{��9�~T���3�wm���E�K��}7��6�
�N3������5^^�j.�E#u�E3	r�j٨�Dv�{�P�zU���_����C:�:zuM/<�ldL�]����=��;Ӷ9&/@b������Xѓ��L&�[)�#�3�S(͚*�"@D���%��ݥP����G:[�*4|�ne��!ך�Q��P�&���^~f��h��u+����
9�B�5#a�l���<3��A����������K�N[ ߓZ?���=��,�5��J5_X�+<g��TydfM����O�SK���|+�I���hӲ�$!�#��SDQ,9H��GK����F\s�	����М&�p���a��'G~&�N�Hҧ҃W��F�qx�5��;����t�g@:&K��37������dBنg��H����1��6TP���yꝀ�N>[[].�c�������~l�~4ȟkL"7(	�����<CF�u�k&�8��y}�]��y�s/�ٙsk��1��������]DsXV��ǼD���n����e3�@
;�0/�j��]вM.��/���diH�Cԏ{������\倊�����aZOz��s���J�lZ�qiP�����N�w������w%�Jp��y�p�؊o�B��eQ�S�Q�O��#�:��4�@m�,��o}�R6����:�f$2l���|��x:�PU�6�Q�3�xIdsX�Qs���z(������c�=\�w~�E�tr���Z��l���йyD��c`jQ
�~�/H0���o� ��b:���#1�C�r8CF�`�e�D2H(>Vv$:��x\�*��D����լܢσ��N	*`=<l��t��}AS���%6e�j�>บ��U���u����b!$8������r���?aB���T�c>)ό�?� (� �A/$N��,�P�Pf�aZ�Yy�q}�aW�:�MD��O-�t�I�3n��(AZjw�-C�5���9Hf��_%`v��Q�4�5^�8i��.�v�oI��x/��]��c��ݿ�G	ĭ	Y�g�&��c������3���Ur���w:�K��x���a.�ʴV��J��*���/ul,xEt�����b����V���I��"�/�T����@�PUzP���{����C�4 �?��ek�a��	!��X$�>/d3{ �X�9F��D�`�搃lr�v��b�TK���q�R��?T�y���v����S�դ\-���1)���iw�(�����w�8��G?f��.�o��3�1�r�k�x���6̟{T���0%��!�o��]�Xxe<�.~�y�s�H	���%��t�胐�P���nk����M���7}�hB�'Q?�Ü���1W��@����s� G���Ο]Xm΅1xs�����[�FS��'���T2�B��֒~V?Ir�eE��W�����Q��}��7��}�]*�%�5�r�,�@^b	AP^,�%�P/2�S���?`u���h��;�
��_z���ǒy�C���C�~��P���Q�"[RX�,��]\�yQf_���'s���/���>�TTL��|�ZE�c�#��&q�����D���M����_6�l�&�X�P��ݪ����U�� �	Ñ�-�-"��h�5x�9�'؏9A��$�C�S��O�ZBjl�2��1F.mZM���S�ğÖi�SHP��}6pOk��$��9u��,���O�\6�P���̖�R�~��	iX!h��b<>�Gz'�3���������j\$3n�6��:4��b � șY<H�"R�E
���p2�ڔ�"d��|l���˻v���v��kv������4��'W��vI,���jDp~�62]������̠;߇�E�?�y�;���F>�r��j�xܹ���w"�$/�/�i�K	1��d}��қ�Ȓy�ҷ������Q��5|�!��y�/k�f���Μ�ئ�����G6x|�Sf7��uzt���rm&Q�L2��:��0�����嫼�ȿ�Fc��_��a�]>qV������fm��P����/�3��X�a'����9
��q��j�YUq�,]��]+Q�l�:���c��lO�_ǋi�L��I�6���m�+��}T_�M�gn��fE�]��v�ұ6�W���̜\K���mY��H脹��޽�$��P^\���W��h%>T�U��6�h�u��C��AS�����1r���%�tȕr�B;Ck��J3!��H�A��|%�ٚ@�O�(H����8��k��ԃ
�Lǅ���y����:�+~p���m���u辰O������7)��OU"�'e�z�+VG��٥S)yp^F+�V*G�����pX¨>BP%;�KO�N���X�m4�y�J��I��4�&����lv��3��k��B�U������8{����\�v̎���Ε�.�a�HwxǊFy���'w�PI�$L������]�C��fֈ���r:�k¤��B�ЂH�l�=��fR���3�w ��BӋ��� �'�o{oz��@�����:-Hvc�#��=��V)�u,�T.�����B-��'�=��x��z��+|P�q0|8
wS��)]G1c���]�w(��<x �*!��8�>���~�����������e��6BD,F�������cв�k!�E=x�]痛��z+i�2ߑũ�K6�1L��J��>�����Iê�W�-¢�
�ġ4��V	{�t�%��6#���T��NaBې��~����@f������>��|�	���2Da+��ɰ]�� V�H �G�H��s�����D;�;v�#�S׊�
�J�کr�LI�B0��V�<�r:��";�S7h��zij<	e��+`7�ZWPʕ3�H{�		�``��œ�L�M���E߾V��9�� ������m�Ypƌ��d�;F��JRԱ�.�� ���Nc� ���w��y�x� k��J�|������#�3Ⱦ�#(�4Iʀ)���5���)��;X[�p���~2�x<�)�>�J�m��!�%�qӔ��8���ণ�����PE%/�ۢ6Y˷*�Ʈ���� �6�ɣ�3�rĜ�|�~��z+��'�$Od����rb��Z?R�����F`N��c�9�c�� ���&��>k�(8Ŋcc �'{����9[�ʫ�o���%>Æ/�/��dOKg��$����������'q���t���x��^e
��fN@7<���;��T��wJړ��W�
�F����X���\\[Q����Ӛ�}�ӂ��?{X�ڼ;B���+�c����V����g�D����ZGd��!�c��*���ӏP��[]x]���L��^Ϻ��t��6\�7���9������ȋ�29V���{����TĲ^�j�љJ��XM��x�m5���}��I5&N�m�E,��@2��1�F���X��:Y�#.T�q���2E�e.�YJ'�,�	�W˟���s���=���2�FP�@x�16�m{��3���i�y�d����Ȥ�η��K>ί�4Z����a���Jwx���ݗ�~p�A�HI�58����#@VHA�Y����ͨŧn����6����a�-&3��ϊ�\�mt ���lU���3��Z�{a�%I�j�4 �	ś��s��!�B#
�{n�:�D����5{�$D�ǖm`><B�b�� �ꔾ�'5�T��cV��:S���;�CtK�:i�e׶�nπy	����v�ſ��!B�w�MR��c�!q�p������#�Lд#f�^ߴ�Σ�q�&}M�{M�.#]�C\5!��֡��/��㐜|<g\Ro�ӥ���Vst龪�� �W���Nd�F�o �~�6��
��_m�͘%�P?&E�������e��A���}��ix�D�y��ݢ����j��8r@�Ԫ����h�b"[�zB	z:�a<2�'Q�����m�u��~�!`� ܚ���A|qP(�Q��)��-���:IhK�s1�|�� [�N� �-?�\L��m��[�ői���ٔ�xѻ�݀ؽI$-�N<��\~ ���jKz�7Rٷ��T	� �Y;���P��6Nߍ����R�l�*Rl�������"�?�����Sih�L�}b(��B�Ky��zӀ�\�͖n����<[WUB�� 1�Q]�/'�J�I�\V���1�`zxI��L"�G}�k��V�^�7�9`ǽ3���+E������\۲�뉳�O2�q�J|��p�T����#L�qd9����Q�ݖ/����x�{ڟ%n?0��2�G��`������X��Z3��\n:#����g�z�c$9�� _d����i?�B���:Ot /�>)���˷��[����o^��MǹD瓀�X�G��L�yLw�*�^�@6�c8���!��,��%�>\�������vt��\UҐ��[6�d�t��?���e�S�1��֤ dC#�k����VK��DC9�����s��'����2nܭv�8�Nf�)^Rߊ�� ,c��MuX>[�oLu'**����ɘ��a��]}8��P#�9�.e�y���ә_�,���m �>e�Bn�˭'ye�I����@K�eȿ�;���^o�J5�������T9�e B��F[0�D�.�ų�P.��p/}힊a}(d_�' �)���$:��}�*��8�Ɓy���tI���t	/O,�t&�fC�f���ӣH��'\����@!/
�p�5��m'���G�m?7�����\^��9?�h���-�r��<�"i~^�C�:|9�.�ݒm6a7�"���Zϭ��̬��  ��h8��!^\�	��	'����w7+^��$�]���Ԣ����ҝ:_C��D܋���g}YRp�?Ǉ�^&(�nh(�U���/�ˤ�G�3��~~,��Ơ�2�Յ��9 R�\���A����4+ O|'��(���,�G2=1m�\,f�%�?�	�ݬճ��{9�Ʋ)��F���>�������<��4`W�K p+Z5�|u�;��������S�� -T~�1����˛&����%��c֣)���'��G%���O5*Q7p�P4�.I꾯)<�BZWk3^�g9�T#P�����܉�Y��Ӓ�p@
��F0[D�g���T�#�8������V�Ѡ�q/Y�@���M�|s>>M����"�r}Ov6�X�L��]l��ٷٯKR�9&S��]���H-Y��~�%3���F�Be���1!�/E���c�^���Q�����쀓�O�ٳ ��v\�~vJ��U��0faݿ���zq�ZU�r��z_N��|䗬��]q�ef(!~��Z��Sn�T"7��7�$-8˺�	�G)��m�ㄳ	�8�R���׉QY�3p�O?���U���[U
����4�Q/�t��#�r]����s��3��T9�{��Naxp���р�ad����o�$U�R��(@LZ��� �%��x�0
�+��(�aӺd����Ӕz�M�W�^3����ʮ��G�R�S�l�s�8�M��G�}�Jj&��p	�J\��l�q^�����`����l�/M�+��A��\�R�I醚�=k0�>��KQ����X}i�2_�t9$V̝����'B������*"������QΝ���x?�ˤ����n��EW�T�V1y��[�t%sM�}��\���أdvv� �ސ�Ie���l��
=ȿ0g�x��-PW����|{��#��G���f�xRz��1� #��,6��-E*������	�	��-�!�G;��#��,�+phO`$� �z�i"_2W�K�&e��2��ߡѨ�˦��Ւ��;�,��O�9Z����d��Kx�����0�T��,j�ڠF�kSфC��4ʈ@}ˡ�
�k�ۆ�#."ԣ�1���x��q $�h��ĵ��>�i?�{���_>���=-�`��\l���K���ᑪW �����߼u�!6��h�e8����MO�I�C��[�ra-XNH�<�	��������'v��I잰����,�E��`�E�g����n/�����`�18�>�4GK�ֺR��B)�0 �"䮇pk-�����J -7G�.�Qy�.{զݶ<�d���Þ������].�):�#b9wR�d��^�����4~�2�~��r�T��.�dU�U�l��Ҭ�)��
Ap��]��tbl`u<���)D�<eR���>�ϊ�o?�Ejivn�M���	�]!Wm<��W!�q�@^�09wʦ�*qk��u+z�Kf�H|~����x7.��E�V�����¥:8��q�[P/ә1s��~����IG&�e��X�7	�Z,��Kςv%��[у-O�eULX�i>������o_�E���m������*	IV��}c����?�
��A�8i��N�Gw�+����WM���Z�#���r��:T��A�o��y'�Q�L�y2��?���7'�)�&,�Z�܋�N���>��h����Aruwt��S�f����\��@Pcj"�V���|:FS�����g7oB�#���,����2��!�Y��v�rM�=S�śR$�����󌎢�&1����KKb�w�s��)E
Qv��<���Ϛ�{�H�Q�?1^a��M�̸H�D�mE�����4��#�K�cPJ���C�G��p�ӟ���iA��ڻSG�qN��k|�ZF���Q������Q�.t��y�����Dq�>�c8�4D�߄(�"I��f)z/������[T[�����K��lw���h�ۈk���r��ѓ��\#ȥk��'�[}�m\C(	�F��2e����4$\�Щ�:#[�n�����}��R$K�[XB��"�$��o�6�UmT��9�r��Z��|�5ӔOGus9�@\�q�l�{�k�f�d*ʪ�@wx{�5N@
GU:�ORٳ�<��e[� %y�t(z��
�l�c��a��唜m�%�H���xym�hb�1���9	���տ�M����P�	ĕ���֮��̤��,��3�_b�qjJ��v�.hE���bzڴ|�ׄ�������d�yZ_)Ӏ{��S�����e���3s:1