��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����0� ����遼�6������"���#�{A���'j�Qj} �}xT	g��F����a��f��洜K%g==�Z���L1������bG����XB�k6T��w+F��3r1#�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^0�"�46Oe���ӕn�K�.�"C(%W�F;c�s|[iMH���1`���TSy��Y�:�c������s���B��)K�����6�K�����=*�;�cWY$�t��;>����~��-����i`���㊢��B�r~L�����1�1�&FR�M�ֽ�����Z� ]�ŏ.B�_`�N"��=���/s��Z�Ĉ�����b`�e��b��S��/���Q�sp3P����/Z��/[�J�h���X'�[h�֯�+���U�cIDy]�z��vMU����~���x�.�+��[i�S�<��ȋW�|H
U�˖fcN�s�K�qU@��=F�"��{�V$�M�*a0��mKo�|�oN�A��yeB2@tt7����&�]Y�sr2�Iц͎sK��x��:V>>�ʬ�V��o�\?)F����\��6��H����)2��	`�[��q�`��UV��(k�^�~��^�+8����Csi��]I5�c���W�-���nN-u�.T�f L���;j�K0����)��
?�����,�c�f���.�_���U�0�}G�0<��.��O�g�(PF�Wi�r	o��
�9��ϥG2}3	�nN�]C�����ԍ��F��)��OZ^;)�.o2/�W��-E��/��c?��n8� x�N&�-Vm�_�nH[�B����&�4�跺�A�H�~����Y������҄��ӈ �mkP�Zql�wb�c@�[�Y�Ф�s�Y�Y�R�� ��ޔ���ʷ�����<I�0AJ�>{5
��]*��[h"n�����\�f��Tʻ��4/q�o"$#7�="ߜ(L�zV5�KYf+
=�Gk�v�L�gwYMY���b�׸�;/�g��E})�3h`B������ٝ	v��$s�\�������e�������8�����9��"�r$z�g�^y��:CY^{�H��ۤ��(�����!s��+b�qO޳����l�=�O�f�6j����VµOmý�#h��x��#~���,�}�NUܺg�n������<At*���͜�:�#[�������Ǚ�l��լF���G:�!bb%t8O�%��ɺ�����Rv��*HQɀW�#��MhBٌ�$ 7i
h�WF��0��@�㐢���ӻ*#|�k*&p��N�2~I�ݐ����?�%��)4B�����+���_�ԭ0 d$K	 �$�������j�j��!�O�;{-8��Vp�5���\����3+�¨�1{�T�Ӝ
v.��J$�d�ǯ��>H28-�i�C�⡔�����ˍ󬄍;�a�	I74��y-	5Ƕqze6��/��9[��`�ŀG�M�)�-�
��?&hXq`���e���	�s�)J���14�w���.�=
s�����l��<�Qh׳L\W���޵{,zO����0Ѣj����0م&��KS
XJU�.�s�� (�%uH�:~`�|����E��Q1p2�!	��.�����G�����lŕ��8��g��vd}S����^1�쑜TN���妄��i!��(�Õ������'(/Ձ����$��f�K�&��gJG�|f4����Go��u��Դ[�6I�j\�@�h2�2Q@нgx�`|V��5M���[áM�@��Q�Q�b@�6L�;̜m����D�3�]�E;���z�fC�x��#D��z>��;.3j�����\�[5xJaX����h�%M�)uŲ2��p-��^�B�T#1�����,�XXo�����^?�OvE��M4��字�B��h#,�[�m�P�R�[���ƕ�K�!�)���B��x���,Q..W�PM#AW#5�������d�P��1�C��Qn����'�=��]�섞����7����չ�V�y�>*ev���2�������C��G�U�x���i˹����
Yr.]�$�=|�ӓrF��f�\���_����d�1����^7�"�G:�^[������A�������<�4r.z������C�����@�T*������/����͢����̼|-�h(�u��I2�K�b�[��ۺ���Y�HtEF��S�mv�h��{�(�!G-����܅>m�&�B��X�E���u�S�$�>:�k�d�~��j��j�J�LB�iASL-�PےX��?̎�/��ttx��� ����a�J��4'HW x��*�I�X 4z{��L��{uZ�b�~�it�-%l3���kC��C�2���8�V�2�&y)��tHE���j�ȿ]���0�{!neF���=�Oԕ^��%4���dd�g�(�+�QB;k��ޯ�z#U���Bi�x�򘏻W����w��y <�0U/5���{�5(���J�km��3B>Hw��{i��?+�����%L���cr��`��skyR�qK��=�݇%��$�>���ͽh�i������ύ�������7�r[>^8�E���pFԑ�of2�sͰqS��/��Rq)}_+?�g!��=�=�쓲_y������R})%jU�ٵ�L�r*�bHX`��{R�]\�O�c����P.2ǽ'��B�=�cq��ک-f���s��	�3c���Zmҍ(��p�x?�|��4[<gE	.h�n�D\j��HI���Yڰ3Vz��v��$#��9���� �e��2��t����k_����k�=D.+]v��B�Cċ�����䲕���I+�����[ ������J��) \��@����2�g���z���f�z&Ô'�hĨ���&"M�C"J
D_z�l[S�Yo8��D�Gn�+���
ԉx*t� �H�k�?�@ґ�D����`��_�k#���W�0��;d���{y�d��;_|�L|�7����ؕ�|7��?��R�%�n.{�+<�0�|bjo�H�EY	w�2���}V��g�Rh������$!�T� f�4�٤*��WH��fm�vZ��'i#��R
�,9m�6� &�ך|�V��gm޴r��}�|P�y��"��FA��Ut�ą�b�&Ԇ�L�˳��h���a���ğ��� ��E�R�e�[��u?�<�4�����?�%�N�8l��F�!��e:T��V�h)�EG�?Dh�e ��)-T�O��M��4�^�yEo��V�"U�c�ql��+�4N4� ���ߴ8����X�5 }��%Rkp�����X��/�,B7=I��F8-R�Ryş�x�4�5�ز��jF!�[� ����|���ci�D�oZ`^��ξ�����,�Ԥ�����]��!�)
�^�A�+Ok�kX���l񴌼�j:%�
�,�_�/��-�#b'|�o���"���.��޶�!�PD���l5}WC:C		^�K��w�������ET�+������(ȲH�0\������dx�A �3�s�-�>���
@�OնS%ȹb|!rKy�UNS�Q�S#tx�6K��VRp"\�d8���2M�B�r��h�����t5/�TW�xE�?�����`GKSr�,l�\< �o�8��0h�����"
gF,�&.�ž6��ݠ�z��H�ߊBٔ�Z���!��T7?@�3�ѭ&�XMKE��=�K�1���.&��
�����F�,B�Mu�˨��N�s��Tf{�"
�۪G��4�R�7��o���.ʃ���� �RNZ0�g��l���15��NjU\�O�j@gW�����Y͟�[��j��ܸb&�]�n|�@��x�{ApI�4��h�7�?�a�=yU�r�_ʴ-Da|^���Eي6DY�&3w���;�D�Qe{V����Lr�3�Re_���7�?�xq_P�wQ'wV�;ң�L[o	�d��^�F�4�/Ĉ�+_ؗb�3
��%u��?�P�Ǳ�t��u���űm;H�����Tr⏬��`��E�k��	.VD��u��y��
f!̢?������7�~璪ܻy�����'S��@�O2?p0k���<���;K��TOt� dFhE� D�b20Y���H��q���������a��>VA��u�H�_�XA��w��:��,s2R5�?��t�n.�n�\�1����[��H�@�Q:y[�uv�ϰ5�KX�Lsۯ��R�.��( d.�0���ͥ$昊;�<�Vw��r>�����~��E�Y=y��4��ş�^.�'4����DQՍK�Eb����`U��`X%�z� �)�H��~gR�F�~o�>�e(�f��D=H6Q�9�U�Tk��l���}���پڠ���4úּ�r��N��,���f�$2쒑rN.F/�,z��|�ʡ>`����3��c���oɁj��Ň��S�.CcKW\�P��!�81������|wI�i���_;+?a��P˴S/��T��ED�2ry)��"� HS���v��I��@A۴��~�fqUm�4 R�'�r[T��NFf�O��N�-�#�T �dvp�l����<�Y�B�/dBWQ�t��#�b9`Nm��x8���h��C���-�F�?�P�ij8g,�{�D��H���R�l]�?��l���7��AA9����2�7�#�~J�c����_j�q��.������v��t����{��O]�){*	�k����>S���A�B�+~���� @S+w�bs���8���"A�m,H��䂌0�&`e`|��p���&|�.',���r�O����'�^n8�qG�v��/@�
<ӭ`�y&����1���9Z�������3K*�8%z/u��y��Qk��̰�ډ�NcQ����
�*�w߇jk6�`�3���-%$m���A*U��K��$W9�b�#Z�Z �/�`YF��5��������2w�Ʉ'�Y�~
?��C�v��:���I#`��c�"�̓e^��K��S���=�g�&o�jNxr��$DO�zƷr,����k����L�w�;.�Pq���1���Őn�`}p����b�8� �8�?y!��s3�ޔ��J�T%-�q3�{�5%��V�ω]��
�[���Ÿ� �_�э�Rc)�u�TM^�>��o5��U, ����UL���R�Q��7
K���� �L�NHσQ[�=/W�@>�g@���JB��H�~v�Y�&�����#8f����Qb�X�7ag�>��?>m����g��u�g��KCz0��-u��9�#<�Rs��ps���s��J~E��<0M���=Kn N��ggPD�A�mi9EE�B���-w�K�"��F8�5��� |������-���G�؉)����7w.3�qQL��S
��e�H��t&�k	� ���T3�Ve��)�	�1��r��Z�6����ա���;n����-�r٪�� �6�����^���A>Ҝ����.T,��QJ
�=Ǟ��=[�fF��� �Ь�r��`Y��T�Z@j�:�v��eH�h�����K6C:⑄2��`�X�}�w閝A&��'VN%���p"��3���(��Pkکû�79דH�#b�B{�]��?O,�xQ��L./�]�m�X����r����\�N�(���(�s""�*)a>^�h|OSH[Oo����0uv��=�zT�F��x���LV ��D�J1`��pK��D��t�r��lO�������5��L�5�\(�f�5"�w^?*��Z�>�g��]W	M�$�����zFO_a?p��J���F�����(�{K�ٯ'�3��wF9_[I�6yػ�|n+�M��=�q�&e��@!������^�7���2���9��ʐK<��'�q:o�Q���n�[���.�؆Z�c�:!�y����<!t���A���DP�w~��8I�C�6���YI:�	�"��A�b\��?�Ҿ6�����y������VR?/j-�b���e.?�-C�O2�ء�,k�!E��e��S�R��kiˎ豌W�N�
�p"�b�5\ai�|fϦ���{�P����(�i�'9��&��!��	97à�4�ऺ��f猛�w pr���e�E�����1��ha�f�(��.sM��K��Kv)կ�1��$�k2蚴;�<f�s���D��w�<@��^�S�$���b+�#�ٛI'�/�+F�'c�QW� ��^M�r޽����xf*e[&y��>"zɚ1�Դ�OKXLϝ����eH?A�����%U]wJ�_J� �evǛ�>ߌ�X ±o!P-�8�k����\<0,唭�Q�}�@/e�Z�Q����MN|��RG�����6�P�����}��7#&_M����,��M6�So��,d��2�g4m�P�d4���鲦��ҧ�e����F�pF��qR�!��?،G�)�l���e�AgZH~�}��-�tLڡEڤ-EM����>�R���/
7�k�ԛ9]�<�(1a�\~����9SZ=�p��!�oS����t��hJ��*�h����$���7�Żw�r�QL�$�!�JŎK�g�Ʉ�}s�!
A�q�*#|��.3vJ_�	Z�'iHE�+�yr��󉊟�}�:ܟB���^r����=����J(��Hv��>����l4����0Dh�o(?�n��#D��8�P߿���9Vm��x��E��g��P�8���I�)��q�&E�c]�f}�G���?il��HT< �Ť[��i�:O����鈑-�D���r��u���2�_L�uU�����ۥ�Tn-e\ �O��܊%�V��|]$-e�����'~�y��z�:���C}D"K�N�����eJ�,���Vfh��SQ�D�C�S���K���Zfٶ��M;�|
�*_���F�Sޛ(�vK"���)�`�-PE%�/���17|!󐺊`.��:7�*'-�|��>O4�1�C(Ԫ�Qc��}FD�l%8zC-{����c�D���\E7<�c���Z��wD�Y_�������p�c�F��/�tP?�eޗ��d��`x�*w��H������k�M�$ׂ�s,N��'e�v��(�=�M�#���ǜb-���O�\!��c��a��4&��6%* {�e�k��]�T�%a�>Χ��>�9��X�=|�A�W\� ؋�P��rapRe\Lik��sL��1�ް,M�C`ѥ�9��U�FT�a�G��f��Kl�)
ʯ=����n�~��l����sP�m�s�k�`Rm������6�9c��XD�E%|��j�Uo�����]�#�,��t/yj%�݌��	n�s�*��v��bo�O�@q9�H�>����k����y�L��@������v?��S�25;S�8��NE�HO���W64���X��jE�[ ��њ�,��?�����r��m�]?{��s](!hޙO�/wƀ�6�1q�t�v��Slĵ�*���>^��c񼾻�<��s���d��G���%�v	r^,�8It����=Gt�p�Ç� ���{ZvA�����ї6��:�oW_��������֩]���exC�8Y0���[��>�&��8f���2�YJ�x�r���M|��Q%��+�]`���T4�*�F��*�WJ"[o�1+c�����t9>Z���׀5��.y���M�,Q�#JM�(��lA�v_�̛v��k@x�H;#;5����V�(�m�� �֩f�-y�sFȆ(���VZ�?u��s�)���1��I��g�e<r�F\C�ܕ�lyBI� ������$1�z��%lZV�;!e:�(���!� ���f�q5����7����hߣB��m\�U�
�M��]�FF�NG�]H0�)����H�U h�A�n���A���k�3[ҏ����|-�\�*Uש�wӉ-+����=��$�M�4n(��%�u�/ �~N�rVl .�G�FI* 3�l�ɥ��ҕ9��\��8R$�ob�y+:�[C�B�6S��|s�66��=��]3mh^��e�n�益Sk�0�� ]a⇰�N��-Ȋ�e�U�yS�n>-|�p�*���S�0����2�S�M�4,x�p����V8e���M�
��0�f�	�P;/�]���ĝ�'��mԻ�E@d��2m��~ҕP�����I�0��xлPe�����;�j-g��aDשSE5�z\�R���߫3}Gw5IU���m�Э������,��Z[wiJ�4:b/SFS�+�(?]DC�E/S^�+Z+�ݚ�h��LLF���*�J~�.����kIZ���gK�t��,Z�2��Q?I�ӓI~s��Zz�V�:����M7�&ױ�t�c�]����h�r_/���M��o}����P��
-@ J\�`�/D�ii#��wF� �W�N����Ć[��#{����k0�L�E�~�֊��M�pM�
����ꜻt?�Α�@ꯡ��3K��e@��:�����w�r�����۠p�j�S>�y�M�I򰐉�M!�e�HB�ViW�i80
=���QEc�E�9�Cp�g��8���g��Jh��!���7�̾ؤ#��oG]�ԓq6M�gmgм:e�*�RH�qZL*�oj�4hnn�䍋H��%�2e�ݗ��P�1�J�kH
�i:gە�桊e��L��C[��E�,��R�+1'�bh���wU��A�h60��D�!��/�*�M��
��W��j>A�[f����)CG�� z��A����`��8��#0����g�i��Ru[HX�&פ/��|��c,8���~�Ɇ����۞�%�s'�_�v��;f��( cn6xo��P���u�^�P��h���L�t�IY�x ���ee'�u?{;%�(t�q�=!�7tj(ۻZUC^%�]��>wi)P���ƃ���y�j��@�1P���G�*��n�a���|��^��ۯ�ɿ?�!f0�� �C4;�$�.
O:)u�q��׍�{D�^}z"s��e��yqCTmJ)
��;t[ۼ�[������j�-K+���ˤ��I��`��[�]��M��[!�b�_�H/b�x��hΨ��C�{��͸��Q>.��b���PPY=�*�����u5$� U���e��P
ooB	y������,�TS� ���R|Xv���󮳱�Z��w�n��c�v�F���:'1�?1)�����)��C�+�!�N�	Ha� ����'���{(F���X�n���A�g5�i�{oT� �j�>��RP��(h��'ә��ǖ/��������nIt��ه�!c�]L2��,?�<�K�&� �=���[�E�FW��`o.�q�R�fGp�m�����b`bV��s� W��Jlx��)�Yp�4B�M��}� 8�7{g$׸Z �QO9sW�5�#�k����G7��.�w��&F}�廛�����J��_��� .2{s�l[���Taiw�H1��VJ>����<l �?���Uˉ� �%�w�3+9A+{��Ρ������]��r�V��nX�ֻ�>��{���0[��^Ҥ��kM��u��(p�V������[�Agޱb�
�m�����D�O��1�	�O[(�T�v��2ɨ�@(@)�K2+��a]�{���7ȍ����Ӝ.�J��[	�����ν���"r�GJ�B�dWt\VV�_�H��ҝ:�H�� � ���T�� /k���w� ��O"�p���X���I%)�ǡ+�qt[� v�@�.�6X��474�(�Q��=ٻ�gi M�ț	��<���׻=�g���z��]u���QB5Il�֏�J~�����9��Fc;���
��߿�+,8b�M�5g�5�am�T��^���Pu{,˭%���+���_����a�d�܎8��탞D���N�)O�
�79|Tvo[�o �f��0���{=ڋ�>���;�b{J#s��}=j҆���x&���(~��<�H�9�����Z6��Lx(Q�z�(���w ��΍�W� |Bsw�8��@����A%$M"Y����W�J��7�qZs��rƼP���<7� m��a��|M�Ұ� *VqGwv	O_<G?��v�ҵO8֖σ�~<���P��3 �w�RC�$�
��lT��8��[�N`eQ�~�/�y�	jX���ɐ�y�2��&OntY�3��j{0�-o�.��;�J�HG��F$�tk3����co)!�^V�h��{�yj��l3ѱ!��a��ξ�w�r,�J�ͅ��]�tkճ~���@�����Q�����闧�����x^��F" ����³c|�ĄXsVs�l)�f�с�-��{����Q��t��E}v+I��Bs��ܚ�E��S��k�Tz���1н�T^G;l`�)q���sҏ@�Q�^r�y�{�#E���ڹj����_�o	��̥C[Z�&Q�5P�|�#w+����AXr6~����n�]���yz��
%�P�/sp�"Ґ�I���	1N�=w�u*���
9p�h�B��H��PJ�n\0��Sf({徖?(�S���wk��Ws �����*�.��Y��u�#����(�VQlQ��S<��w�!~��'h���*�[�>�3`��T�b��F���\@T�&�n�
�<��=q."ҧ8�B�x���Iui�>!G����F��׋0¶Xc�����;�F��=�V��(��K�>�
���� ��Æ��C�U�>uuJ�
����H��ɣW�2��.��l��8�.��+���t���z��0V�P���-�
��	71��nd.��~��3Gq1��rÕ�Z7�M�n�������V�c��!V�' ��0e��RG��$v�mC{}{�Y\vR�^�}���\|��wa*��OpAO�)5uR֧]��C<�Zw�G�MmWӎ(����]�D���Ћ��"�`��.���\��> Yڒ��74�@�ΰyO��	��x�^�4b/c1M��K�F����U������4�.F#�~�p��,���G5�f8�	����?��UǤ=B2��˝G9Ǌ�g�]i�"��9*�,�I��R�{%�7�J{�;QD��Ze��f��g{�N�99Jf,L ?�P1]��AS�3a;w�#.2����+�k'�(���1�H^x�B�S��6��ݚ����Eès�� ��ie��Mp�.&���&��f�OתW��D/�4���MQHa&���*�J�rJ!+��/;��M3��@���r8�w;sE'�:�.4����u�[o�_dPwj���t�p�[P+��A!c.��{64�?�&v�`vTQE*�p��<[���sd���XY�ߗ�ioL%Þ�8�.&�8�r7�;��UJ����aI��1u��5�����3���n�����YG�[�I"�l�=!I�6�{^�Bf2�~��nu�l~~�GOu��JHdOR�c.�(�T���R�~x�� �f�g;?�h�jP��Yf���K:֥K��&&zF�222i��j=����������W�r¶���v`5j�L�֜x}N�F:��M"�|�J Lbf�եrT�v��]wR�U�#���iQ�{�38�K��.����e�硶�YM���\��v(��*y���=���Rq�Ѐҵ�����,��hZp���<�ェ�Z�i��))u�kUxnx�d�%���)Yg#ub�2IMȬ�Tk%�R�4�6.n>}�do��:X��6�),��)�$@�p�܄��;w�s��n��F�
ɚM�/VlsnI5�>��H�k�n��x߃�1��b� �� �3C�|8�Н�!w��$�$F��U��q ��#y��dݝ���
�?�t���c�{���o�:��0<&F쉒�d�OR[���٨�wu҅��W��I�H]�~��f Ps�Fo�"�%��� ��p��؉�D+.�[�&�m@Z��7�}߫c~���6��7�q�ݻ��Н;����Tj!^�&�������[��2�;WIsFc9d�s@M���x�(m�3 k��N�r��p�Eߧ��`��Y1�w`7a'���������$���4Q���g�<h o+(vu�>�Rk0'&`�,�(-��@�$dQ�7�dK)m�:#�Rp�\��F`��2:��6~�սD4DI=/��S�gb�s� )_�L`��d� �ňv��u���[x���v��WV%L���Z���Y�&�n���?�V �2xN���d|
�U���?\�ej4��Z�����Yjgԉ��!a�s�[�:o��o��<Ҹ��B�B��Y�4�E�G櫆n�70�ɒ0�[V��.���h��>�������({w)Z���|�
K֌��AD��"�r�<4s��"d@�v>ش]I�Ղ�JBS1+ݧ#�(��p���m��~�t;����8,�Z��ٙ���t{�G�Q�"U�론�<ӫ��F�'�MP�L�0���'&�F�����g�e��c�w��W���áVq�&۽���b�4���G��������z���uz*� �[��k5�@�a1��L��{�ҳ(�u5���>�Ȉ�i���ܑL�x=�C�1=�x�X�D������F��i�@P+|U>�B�F�>���:��b����E�L��VFlqDb�E���c�+�'t�=٤8w�w�N�$�@Q�K4�`�uҞ��k��W�w��4v���w<��g6	LN�T�]GҤ<�OR��!�]�:�˄I� lΘ����]>�	³R�l`��@��ߍ���q������j�"��i��C��#� אE#�`!N����Y[K��.��VϠ�t���x�{D���*�U�7�Ym[r߮���$�g�> ؁�b%���J�a) rI�r�{
(�+AI�Tk ��Z4�*��T'���Ǖ��DV���2�s�S��5[����W�@�Y�+��}�h�Ӓ�"�ϑC�-/m�c*V6�JUk�5ɾ-�.yL:`�� �:v3�!���m���-V�:��f_��ޏ
K�g8�f�m�m�qo���v%��1j=�x���>}�)��P{YZ�g���cY��DhdR�1��
<"�8�S#���C�U��>)䇖V s�'��{%�m�aK �>��j�m��o!�]���sWᑷ�7��2C�&�7�I� �Cտn)ǉ�bp
��B��&��Z��+�z��bg#7��4��Z$���so^� x����Ϸ-;8[�c��p+N��l���jx���;Z��|��/X�uq��F�R��3���D���@ILe�K��H͓Rp���;u*L˕�̵ p�}��$�����!��	 n�p5�����p�ض.�P��fuF����� 	m]�� �ﲹ��ň"b�p~�1�)8Ȋ��g��A��9�|3[�lE� ���5#�Lk���y7���B�X�}��qA.���å-��_B�����˔'!A4��̪��":.cF��-2��oZ1��}�&��a`��M��5�O0Xգ�a>@;���C��9�����'t$��<����E�`��2���aF�_�SA2u��0s���Ѽ􅗛�נ�n��ʛ�P�F:*F��GĦrv�*#���ʽ�Y��bP���>���b������ЪM#,K��1�C�	}Z��T�O<�[�~�8��{���LG)� ��)n����3R�|G�"ˋ�����Yڍ��o] ������L��G�u���>�}����=������4/oz�eO�a����0�C:��g��چ@���)�8��r�ƒ���!l�im���J�vp�|�ef�(#t�ׅ>�H�)g}O���Jh�6b;�!iM,��������B��� 6�f摙ͫf�o��O�(�<�TK2/s{�T�а��:�l�Ӿ=�SS����P4|�hTZ��#q8(sO\Uz/ALUwr"�H~p�(C���7�!s^�����x�\p�j�J�a��u��������'�����1�Ԝ��A��Dk��Qڗ�r�S�A��1��[�!�� �@����n���%��-H�?�L�ۥy�],�^e}�x䍅fr9� �f�Υ�LQ<D��#�P�[��i�>F�w�2�VO�o��fk�|��^������r���F#�������9���G�z�{]�͂��K�^����f����g�m8#8nl���y��MXt�:`��.,��,����T	�/��`�6�ȳ?��L#J�l����*�2�4��/r�U�5u�nL�5Č�	�<�>�Y�˒�\�D��wϥ�ȸLS�$��'�R���T(�G=|��dx�+rM�-�~
g�=�	�ʔx� �|�߼�4�a䜦�pQ��>�� <`;��Z��u�BуӘE�$�C�R��������c��8�~�7��p�f��8i�%�������ZT�	`�r���4��V�bOQ��:���b�H�-^	
H��Ebe|<n�\�TﶊK�>�yk� �ac�`����h�	F��^��}6`���x��?��\��ۏb�q�U�����T�n�d����fz�<�dr�;U��Bl�&7b�π^��JM4փ�M�̳�H}���:R�z�Θ�y�b�' ��~��7Us�q���T��^k��+���Yr����-*]��9*����t$4ڊ�3�uM6q?#�^oEΥ�>���.&�
<�5��K)�t��i�FQ�n؛jU8�w>�T�dJ�Y���3��] @J�W�o�1�	*he���]m��ƛY���]K�A�.[���S���& D�/:pu<%Qu#Һ".��K�
���e��/'s%�5�pwƒ@F��#�T������3G,Ѕ*�e�  ��3���&�G9�P9��4V���8^�SN�:��Ô��i|fe�#K��!��|���ĩ� ��Sֹ�[�Kd���������E$о"�N+\wN̶2l�CG �H�>&�3�뱚����1R�a�����`��j4�2�X|�쬥[�9 qsj�R	,q;~;-7O����Y�5/I`R�1G��v��v��LnW��2{yu�k�ՠka7ͦ����-��\i�$2�nX�a'�Ӯ��r+��VY�_b!����Q�օZ�]ϟ	��̰2��]W���:��[�m�hu��B�����s��"-�KOS���]�{��fp�Y�2�Xx%�1�b�r+�����k'�.�������Ѳ��S���f�}��)�`�SKnj悆=\���*G���'�(h�DjG�ߖ�7LZ8�
�j��������p�(�<�ʾ���{�WDo�&ȼ���XÁ�$csZ]� '�%���z ~���Q����;��f�2�¡��	`m�d�8��a��t� ��ñ����w��N�b,U9{��KS�)�I��'��s�o�uay��db�h�T9����̗v��)��cq���!����o�x�U�����й=4|�<!�R��n���^����a>�0�\�v�il��wP��lᦸl��Ķ����9?���w7a��S
3����k�G��U�F��P���7(��ȹ�2���+Tz�;�x��=`16E�NǗ$j�n3�i�/���̔}���h�3xpD��XJ�\�> �P����@�e��|��FtHO$�)���a�V�3��
m�(� ��/A�ǧo�A��('�yMB���-9\qNƗбͥ���{�����y�[>w�GΑ���qs���Vq�Kz,3yV��{�A�/j� r�HeY��a"�	�Y:B���;��r���@��C�CFAW����%#&g��}|n�b7���kd�ů�QCF��Q/�ӻ��\�grF�)�[Ɍy��Byy�"?���e'IkԔ�
9�{m�('�GG�q$�@����gf�b�����u�2�ʞ.N�/6c��^�k�B5#ލ2'"<[��|�B���N�%#�����Z&u�ݛ��2E��p��n�[���]���C?q����'��(��q?� ��h��F��P�R�āhF&��A���\.�`� ��^�d�e�ZLkY��Owu<W��2��)+uWe��m�%���n*4vj��>w��]<˜�����<\J�%�]g��Z4��O�"��\��֊�ǀC� +tZ��a}=�!��[��\4ĤQ[�zm�����ow7���آJ�C�����I����qZ"�,Xv�! �L�)�̝'[�5V��.��a�c�.:�kz��!���Y���9BFV�o��� G��)!U�Y�ՌA�p>X����a��"�7�^���a��b!��,��O���L`I��<��P��o"[_r�$o����6B�r��>��ӈFB�,�Ccv���:��xf9Ȫ)[�O�9�8��Bf����g�_|U���zA����I�H�\Oo�!�2��D�#Ċ���n�[_',��3U���b@��D6H�şCK��>�p�E�p?6.�V�a��VcxH�@Aǝm��o���V��d)��c�Lk>h��q.ʹN���UO�'�V#!\��G���~Nm�':"�����?$���[�e�<���3��%�e>��u����B�����( �ߖ|�?-@�*�G�=�1ؒ����tYzl����x�H��Qu�h�H��_�%�C�Y�� ��U��<��y-d�����:
�ӔWnX+-q���6/�}2�oIX�<��U���q�/��׬�����i�#U��Ѥc�a�2��9��M%.�j�5���˽i�]r��F��DJd�\0��X`1��C��~�7�g2��p� �6�u���ˌ����V�nT5��U�aǓ���n�$� -���+%�?ݐ�z�����բr����^�u���k7�j,���ť��Q��Q}P���R{�=#/�����׆D_�q; p�/IU�J�+�������x�dVju��x�:�Apw4	~��w�R�T�'�L X"���ר] �/���(�"��e��-��̿�զz���Q$�7MT����p��
y0G�Cq��qd�ƨ�ޙ��@i>�j��/m����9��_�����(�:i戢�|�V���x����)Ac��#6*rKq�{�2�r��kv�a2�Ћ��W0���3ٌ_n��Д w����+ �5Д��c��Їw޵�	�R)&�`A?��Ɵ��T26�mhY��a�F�`�6�#�c�ʐ�H2�F�,��V��&xt�>"GL�m�D%j��,��K�v�"=~g���ȟ����}��B�H�فrR�F���=�a:�� ao>SW��퓘h/���4e�PҶ���~i�e�<V	^�<�r��M�U�Xp|��	?Ǣ
fZ�zB}�V�r��I�ihг���^�1=m��C}��~ȲdP��H�A"���=xA��v9��c�]��AAG0Q)N�$b�����)1-O�N=���Y������L�=�$yz �w�J^ׂ�qz���zf.�#�����X�10�%g�f�������y�_=��>V�����/���i:�H{�HM��BlJ_�
	"��nu�|�h��C��>�s`E�t���m�R�0�������{r�a�~�1V����d��%��4=+Ӿ9�{��� �ɬA8�2�[x�g~G^1`�N(��~���!$����.HE}�^6���Xr4��<�}r�_͕$p/}v$���a-�=p�N��M�L�*Јe�X�Պm�e��Jܓ 3 �{?�C�
�����&��|)�e(��_q��1�G}))����5Z׀�ټt���Bp�s���{65�+\�>p/���.
��j�3Qci�a��[5}�B+3�pPg
�IHCpJ�=R� ��5��aV�V�[yz~��5ܖg[�@���'���*9;�X�F$;�5�r-��]�U2(a�"���ur��\�+��%9o��L�/?U�ٓ��Ր��E�Ӭ���j�J���'�t��Өn���U�z.gX.h-vDޟnd��9���O�L�O+���-{�;N=Uԃ}�!7+U���㬠k�1�@צ��R4�@3"�^`\aL�RJ�F��[q���g)�$_WSp��|	�cT( ,	�5��qm�Y9C2���;7��bO�0��5��������i���/�rV�\p���"WlJQoP�'��/5ǭ��۪{���� �zL���d>���� �>`��[�S8��xs�BL�=�N����#�����淪8�������4�S�d�G�H%$�m&|_�Ŗp���:B�@�)w���f�c��&�vm�\z�s��5��4�W��rڵ怆������2;l�@�NW8 ��6�����І��'+�������Ī.@dڑ��$�Gl�����;i�D�.�S���&�w�07I��9��o�7�<�a�n�N��N=?-o�/3A�)�r�b�,��kd���T!��a!���l���(�Nv�aFs(,����B:g�u �5�V��#X�?"h�
Ƭj-S���D��6n����C���M��D�6��N>��,�j�=~(�`�oH� �3J�{��DC��$'U� ޑI*�oWUG���~^w�gM,�
��	I����v%1Vpv�z 5i?�M�2oi�:R���+(��)x���2�����;/
����:Uk�)N��~^T۞R�!	��	���kE��Ln�A��AZ�n�ã��:��Xv/8�����a��߾�ã��Y��c�1�>�ã7�!6��Ѹ"'~ �WT���Pc �aT4�zK�I[��wtk�iv�:xU|Io�1��E��I��%孷?�_bAz,@��u},�0�R�b9���b��3�
���/�H1�T�����a��a�����kÔ�Yń����iM�t땩��۩���cok���l���N�c_��s�g��c�P���Xg)'H㕅�� ��,�97IqY��[Q�tK$_&��;��́�W�!���4O?��Џz�~PK>V����\X_�[nF�$w��ѳg�2J��z���}�,qt�є���qZs�6DB��"�	�됛�Ysn7U��g�d��.	8Pg[<����^.#H*��L�	6-�Ƨ��O���l��~ݎ�IGÖ|��!����֦0�-R�F���)�%Q$��+��?��'�ڵ+���i��7pv�A��vk��c'�Y�!��&�׼����`Zt�X�7zRVTN@vlAP*���
������ �ZK*S��(?27��#0 bH&�����K����l���#�Q�9D@Cq\�HK�����r�+8楘����zr��`A�;ߕ�_7�9z_�8�,����b��+�Z])fglx�B3��;E	�y��.�G5�cp>u�������-dDX2y�ħs�h���(�?w��]���R՚�����Q%��Eʣ�M��*��׵ѕX��<�$��$)���~/���jT�"F�7��E�j!���ؐ��(�E�P���ٓ�w�[�,j�W�粑8�#��O���=�CWG�\�?�ˠP�/b�-��v�Tx�c4��sTp�@�x_�\;�>C���,�+�e��y��Ӆ��Z�T�̈́���}gx�FL% t���M�:Q�|�
G�����g˥bv�H��v6[4�s]�\��ڕ�>�jDl7Ft�|�Hs�r@�u��)vl�5Ac~��W��9y2�-�gf/mc�q�,;���y=CbT�̕*����_��"����P�Ok���Z��t3�T�,�K����
�9�ٻ�@�"���������A��Eўܢ����1*�J��EWQ��	����Z�aӦ��:dL;��2��1�r�ٓ�VT*�J"��7.��/7>g��2:�v�0�㍻�w�*uh�w��xѹ����r��x�K�k�O��FY�&�?������2�,�Z��
kDd�O��"�h3�˟K�YP����c�O��&<�޹ūCL:��*ΐ7��`f�*=U�Q����x�b�/���a��]�����M�'���������!�����V�<�9���+��y8���ç.5�����$�F��P�\���B���1I³>��,r���	1,u����.)/t�E���j�������e�� =�w�Kh����>Ԛ_]��&}b4�� W��4�\E9��@���z� 5����k�O� rFX�l�