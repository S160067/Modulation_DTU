��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����0� ����遼�6������"���#�{A���'j�Qj} �}xT	g��F����a��f��洜K%g==�Z���L1������bG����XB�k6T��w+F��3r1#�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�A���0>�kz��/ �_M��<-�[a�%�����'(�S��jS_�,��8��T�.B߫C|��N�(ݝ_l0fS!��mYԥQ��DF�S;���h/��9mϓo��ޗ�������t�a�L����H���%�Rqp���a3J���Jpچ�
7d`��� �n%�4lP�*M+6I����uc#�3��;�^���X^�=#RB�Lz-�Hl���>(@�A�1D\~vg\��f5L!��+�[��a;�xl�]΋����4�dn�g�$�5(>���|����B�&��cY�/�8��
�E�̾��Lժ�3�5?���q�W��"�0���WBVӮf��	�Ʒ�|i����ܞ���_bX���1:��#�%�M�����d2G����j���℃��ύ����D�^T��;���a�r����;��u�*J��]��4�[�� Yi�1s,rS1��d�Y岌Y�i�mѦ#.TC��xvc���	�x��$Qe��	�>����=*9�W�؜%��úZ����--��:�N�y�9��qҶ\J�H�.�v�Zc�C/�7		RSUq�}���zV�@�= ��O6�-=�뫼�^�XJ�\N����w;Ԭ����7���o�Š��~�4�s�����B�s��#���`!�j�w�>|k�#}b�x�<N��a֒q�����!�΄�T?g�8���T�5�2��h�N~pE�
�o֙�¤=���F��X�T B�6w4�X�V�)�������JL׊�}¡�Mx����Q��h�GR��'���8�,�N�<2�,�G[��Q�>��])�tE_sw�G��P˕Rε|����[s,8&�����O中�6����L�<R�r�^��mΊ~�c�@i�{�O���#ƥ2�ވ�L�8B[���}�s1a1��P!�m���$4���!V����b���  9��� �Χ6.�<��ZL�2�S�f�,u$����oEď�;ф��R@����^�E*Dp�b��N�ߊ|0�7��n�������O^,�d��:�q/����A�"}u��w}KU�+�k?�>��༫���~@���[_z��q]�]����K��qK��,u�_UĽ�G{�C�&h�=cFEo���e��=`���=�	ۜخ�LI;��L�I�q{�7��`��O90��ѣ2���b
��Β�.#'Y,�$7��2I��Q�mZ��p�x3�)�)��0���z�Sk��Ib���C���LX@�u[D{��L5�O��������p����uP}S��i��jb��k�'�dnD.T��PF�V�pχ��~���Z~�Α�M���Q�t�Ib���p|���:/L4�?�[��A��� ^W����Z�8)g�W��������h�YO�+����$��n�DS	�i�5�Yߞ��*V��n�	4~�=�j����]a��@��e�}~gC^��g��h`h�N?�t�c�iB�:�9��q�jw�C��y$8����]�>=-�-qJ.#����h�Y9E>2�lь�MA�z�ΞrŲ�[�`�o|PNc&({�m�9��Yf���Sx�;g�Fw�G�n6�����8.�a%ë��
���Funx>\�;���|$4���-�;`%���˧�/�k�@�y�I\�o7TF�
E��vot�P��a��D^qЮ|�m���c�����aFs�*ze���ey+Y��X�k��hjĚ���l���n��8W�c����z}�}���kZR;Ư���U�1Q�����]{' �Ǩ�5�	���ǣjU���c��:�a�����A��m;a�k/~�D��^��t��=���J�cT�ӋE�6:��+�gdߜ�f:N���ATY������l\;��,�Rޝ��zٽP��d���'߼X����]d/��,?�{JJ�_5��/ԹFf���WGn���dF�3��*�[��fV��M>"n�<)j�Y�b"����d��]\ՙv��A��l4������5����Z͠[�:�.2O��L�����LF��U�����[�Kz���Ҋ�S�޸첡�FK.���iJ~�$��X��$b��#Q���<����n�Gy�TEu�3wNM��"V=�<��<'ǆǃ���F����e���NIY;J"�;1�AsI刨���DN�8��2��:�ZA��e����h;k��\v��-��:҆�K-��/��p�g}�����s�\J������݅�E����ش�esP�����Z�Ȩ9qU��}e��>���~th���~��%��|_ Q,j���g{e���}�sb���
�(mXO����&8����%�6���Cb�/��1zjo,(����ߚȖ�݁*��(�7V�w���Hp��Bo�pI��N]�/A������(z����g���r�o��G�����cta�E��i��G��,.P[�v�z���2Q��gl@]�4j2ç!�I�?�~��ׅK`Ǝ]�z��V`���c��8��i���c��CMZ���K�5��c
�fֱ��߆O�@��Wu�6+{�K�%��`e��Q��f&	��ΜH�in�7e�����=F.As(j�+��ֆ�VW�l��ËƶG��\�Ԭ�t�r���]9~�����R��/��!��H�j޾���]O �4Ew������j3���M~F��M5�MA򊭋���L3�P�LKf3�?~>��c�H��2T=�xI�����}Ys�`���V�n��⛤s!������T ,
�►<��T�9����o��)���Ǯ��
��aN���5�p+kKM�� D����w�$<\�i8�M�*$ ����?%=>�y-G��כ}���X�S��!�Kkq�p�-�$�F:'���L���2��Pf���qEh��Vf��E:�LUj���	@�UI�Kb�1��"��`�fygg*7�/�Mm��B��1�u�gqS�C�wbf�\Xb�P�#$����
^���!(��0��Q��do�������qk8ˠ�\�9U(�j�4�o����uA�J��{r��Bg��2���2'/�<Ȥv�_�?4dLf�&	�{�L�*���_��-Ƙe����)Tt�:|�>-�y��6N��f�` %����M�	GeK/e�ze�e�v񐰊��,		����k����-�����N��O��Ѭ�\C�s��E��!�>�6��L�YfZpW� �j�.OX�S�XllRF���`oQD; �ƫ*�m��7��^�A	jC����"���z� �Óg�~����s��ښYs�T�c2�ь�g h�&��Ľ�[��,�e�z4=�����a���w}�CB�>!T��B����,�Ĳ@C�2<�l�h�v�@2�q�x��Ew.3�Ph��Q���&=�>lm���
�'Q�XZ�ý�����6��>ܻ�a	�m=�O�(Ӡ�څ65�@�ħ���X��us?�SOxA����tH���%O�q��1x�WY&�l
�&��g� t�����r���ŏ��L�*a���P�ZZ����umx�=s�]�m��<�')<�\#�ʦ��~��92���@ahB,XlH)N����
�#���务�F�4u�tZ?��6���P"{k}�$c�J-��>9ڢqz�T�w�{"�� ��P��d���Ys��D~e�Ə5F�0�,��H?�u���1�������6��"mm+^#>�X�4' Rfzz��MP��+M��ϙ�e������'���m��7���ZtG����ay��S��d��pT;,"������Ӑ�Ϲ�U?�m�k�ms��ߙ�3�A�F�$�$��x������W�Z�8'�Ir��k2�TF�u
}}�ky�vZ�D��pH�|q(m�U�����:�ɡ�(a�u��?�O���и����CoG��=�f�`�:�vF��W��,�Į����jƫ?!��P��׷@G'7��D(J�#�����i(�^w�o�Bg2/�?�)�6�������-����S&_��gY�U����-h�P���֯35��W'm�_T�g�����`m�%��W��S]{��e��%�)�C�wF�*�����I�������gE��S�6C�����2Qt���0Z���=`/���b��ڟ�|3 T8}�I���wVmv+�!�-ƣq>w�%���@˰^�,�x�+r@b��g��k��P��)2)'��;z�c�x�"��6�ye���\����+��l� ��s�h��y��k(��$���2�3�e�F��w�B���D��4h�%��q������ggc�g����j�I]���`;R���u�&�Ƴ%��(08�״Υ[µ�T�b~�ד6Mrrl&���3��C_�Y/;I�a����j���ջ4oZ��4J$�[�B�{h��hz������0��D3�\wc��>��p���-��2O��#�߻BS�C�P��}��A��R�	x��}���.}p�,�����5��8C�!g7�랼��`��5��Cy��rC�#C,ކ�n�+z�~cئQ(ر}i�baw�lZ9w�����F��L_oDP\υ)��^ ��o��^�{C�)߸w�p�n��M��?�Y+�����܍�J)�Vs_j!����!K���ڄ]���o;�8���暙��g�c����HMI;MK�j/��L�Y�ٔ[� �@���������	����x�<N��<�=_E��#
_`� gGݜ�+�d<�_�j�����W�E�tP�yp�%1R�*�"6:|	lj�m�d`�o`��rTN?�0N�����.]4�?����'3� z@�(��/\�4��B��0��-4󋏡nʎ:f��?B�`Ȭ������;]�*� �9�D*��ZB���� �&��>^�͸�;؃��HGbn�,z��h:c}Ԭ�u�*�Q�b��3yT��="k)懙����*+���W�a����t.\�zёDrE���b������`�_�'o��'�9��1yJEY$Ml.[G�5o��L�����.ݙ��Ʉ� `�$�@���͞6V6�~�g�E:�A����$�59z�O7vmw&�~[�	�W13����n�;qdǕ]�5L�%��&�Sw%���Q����E�)��mrj�]�ǵ3n֮���l
s��%bi?�J
*ѐ�ONu���}귵���
V�R��p\���K �I���c���D��~��0,�M����e�4�+<Z"	e���ÿF�ԏ����>�j�/u��%;�F�c�n	=�[�Z���hҺ���pʟ4'"��-hQf�$�y5bReT%��?����l��CƇv�z��r����p�x/�����
�j��S!ʇ1�-��l�i$�XϣT��詟1�sU�fq��f���2`s�-���E%C�J�F�]��!��v��f����c7��6@	;�hf��o����� ;���_aKN�](N5r�V�Kk��}��}mȪY��p ����=�kkd���l�GM�Gn�v�z@@���x�iNb�,�Jg\��5W�Ħ{�C�9�pچ$0�p�<;ŀ8��㙁��AP�����A$Kx9�e���-ߵ(f��׶���z|�I�jS �BR	ޭ�9Q�S��'tbJF�m���iJ�)D8�k�}��ͺ��4�O2t��Q���\\�T�T*�<k$ �G��P_��x7�g�0ײ�jˑN�(|�%�y�TD���r�m�U~
�l��j�Gxd�Av]��hP��>�mbb�����_n�6}��6�-�M�qN�K~�=��������J�"Z���X���J{�m
�s�Q	�l�nx��R��pS��@q��+$G���x�Y�E�F��S�Nم@Ҝ0 ��%0>�'`*�����qn�T&���*oN�ql"�c��0���v��k�6N�%��\/��u���]�Z��V�u��\ ��l��o��ݮ	�K ݇g��0j�40@��z�̺����К(}UA��E#o֊��� �g>�Q7�}s��H.7��MipH*��Du�;Nۭ4�G���Wu��q�Q3�;oG�4�|#j6��r����1���;F����]�`u�C[�v:4��vg�MϺ����?�-��vNԢ�4 ����T�&������r*�n�H'�`��0�Αyݻ#�[�X�z�b�˳�a�k����,�Ӂ�����'�n�x���M�;�:�4jԝ�T�+j���c����?$�TA6��n#�8�CYC˙��5���0L������e$Ns�D�?�XmR�4��(��J�h(�7�0ݿT��%�$ZY�3~�UjJ���[�#lyɮ<���Ua��Ԝ[����� rV������	�p%����y��V����]��ZY�և��?V��%�3���jV8�I�7��s:�Y�S��7k�>���ƿ��}E���F��65@2�����!���5c��Z��H���\�=-����Ý�k��v��� uS]i<���NK5��\Ƿ���`�*��ˋ�i��]���$>z��VM�;h`}�a$&cp���ݕ�9o��k����*r>�:��n�ߐ��a��aJk�ŭf�Z1�	:V�n"��`��F�w��,]�g_�m����n��B�B��=�" Kk*�q�CV>��[���)*c��\:֡��Qx"�+���-� t�Wf��� vQ���zd�W7~(c�U܈gۜ&)��p�c<�/!=�QY�u��3��_���ێ���p�>���|M���?���5�8o�w]�*�g���)�)N2a_���e7�	�z��Gݚ	rmA$Z��*�!��v^l�U6ma��r�t+ hF�?�܂��5�T�����>HBQ�� ��$�
'3�B���q����{T
��&_�Ӝv��P�璁%Y��@�+��a%Ӿ��>Ʌ�q_9��l��E� �T�))V�3Jq�]����{�?����������c9r���tփ�PF��G����o..8��ۨ��5�]����M7�-�Q\�Fe������a��
D��.C{�䵯f�s�YPƯ�T���m�.R~9��'}$O�<y�<���-9y��-�Z���+R5T��s��\�ұ�Y���c��!6�����bS'M>;9ؓ��0$nGw�u�)���e駩�6&\�ӹE v���]�LD�s��F��f�tŋ܉�T��r�hp��f���Y~\���Sǰ(0��Ή��R���O�o�.�G�X>��f���֎n�wN������������(_Ӓ��o�d��,ק�ΐP|���X|"�I���N`�
O;��r����}��/�:�"y[������ T:@��%P��p��H��k��k ��e#[Jp���F�>@�L߂�P����s[(��RT"T��23�h�z�Z�Fn/����n�'��/A�[I(-�aj��Y�~����j�f�.R8�
��^f=�Ҭ�{�F�����$mR�R��}�]���QE��q�>�C��Hn��4"��-U���9,�H-� ���>�;G@����Y�Tî(@�=�b�Y[�.F{�9�I����1Ч<�cϛ�uX���>bZK@qW��R�V�*�u�AG(��%W~�8)���`�+�8Q�O� 6�3�:H���?-�_12<"��'� ����Н����'x�0?��ϧB��T�v�B�Gm�VT����ce_'Iy�5Uav������v�~*�~�2��Fr�D��&s\]A�mNaZ깎��n�6$�\�s;���nFx 1*�K)���3���=�a��YS��0�㤃�R/+��>	����0�p�<�"y�����?W9'��-�XF��C30����m0�R5ݘ3�O�xxt���N<�t�ԏ�9">|�5�@��b�
+ÆД_`ŧǨ9��2թ�˸�4;Բ�L%�Z'ʽ��؅C.FcB�vA�!�e�R��鹘ڇP^�n~� D�?b�Uٔ��$�6�bV�@�_��]Í�J��7�w�'QG5�Z�9:�#��$�sTcbO�!=�V����u"�dh�X�&i�d�t�U�Cw��r��eZ��I���ۇ?A�lv3�[���	X����G0a�䇁�����OJC�\��5u������T���ž#]o*��<d��&Ømhb����)'��eZM>���d�#��.o�I���лU�	�'�m�"���fbH����/��qݱ]��'�Վ�X���ĳK�r	$wvW*�o���F)�>f�le�5�-����\M�Ӎ��\|=��RB���7��;+�'���O��:,*����ه���K�Dpѻ�rs���z s
��KU!wq�����'��9>┫�g�`��{	(��7��8SQE��A�{�G�?s��9�pI_|g���71O2Vf�[5)���g�m�?�����3��<=��$��!�u|�-�o�V���k5"��r�q�7۾.O���/����W4����JH���(���b��ޑ�_,r�X�0,t������_�>D��B�X�(D��6���oL�XÖ)�Љͣ(f��4ܱ.���}YHd$���3���B������B0uF��&Y-��Ŝǈ�������J�ʪ�}r�萳aIe��` ��LҬ �*�uZ�?g�be*.&��B$����"���ݝ~-���@�qu�r�. �|aw�d�֢�̉��D��ʮ�?��� ��lu�&[�@ .#�D����oFn��e�RR�D���ʹq��fr<� �+���p��W_�
m�?{��I޳����@����l@Wu\�2���>��3���m�s[������=I(h���P��nB��|4���o�tŴV���޽n���.�&�7=��j�؅��(��������Ow�JI>��R��R�o9��4�{x����󔺿���EW��S\��Ȑ֒zvzj�KEڏ�'��@f�r3�/6@v����O��ڰ/.�(�:�1<�ԕ2&���6���+��hiO��������� ��7�_�hG쏮��iЦ�����\��$�fŘ�:�[����f��A�C����J$LL#�boK�L�8!�"�Xv���[T��ǚ�&ZƁc��8��d���!X�ܗ�PUS h�$�B����+�!?�ӡ�����¥c�����i����ۙ�Ք�q="�\�[[�{I�Bk��>�ߊ4�����sZ�CQwQ����&F�*��ȉ���B̠JEa��+1WO$$]�=�]f�T�9Y���)�=��j�2�y��'l�
4�}�Pv �6�����$u��討�a{�r���,����5��PJ
|����NHGu�+�9�m�y-�K
�dm)�����}J9u����q����J�^�er�^W�@���0D�g�1ލ�흈�P��=�"y�H1�9zz85>�i�fZ7���!�W��I����%�]K��˗���m��ceC<yJb�i�0�,Ez��9"ء�&��N^�UW՘���j���`�ފ��>zQq�H�5��A��q�B,\�x�ì���#q�G�/N-�~WeHR��,������������!b'/�1�������5�^�	r��]�(V�%�	��̝�:#3�eG�V�΄�9��P^9�E)�:���U��뤺a)��R�6;�q���pVћu>	�醙G,z�r壷/!�2 ����jo�zL��	��5�6ħ��
4��7)(����1��YNY�{���T�j�
�#T�W>��},3���NL �k5��m%>kǯ��@t�;xL%�Vd�+�R���̙�(��Pv^�هU�z��e�sѝ`��1I��#eؕjS��@)��z��:����>�
ݧ��4�{�{��O����!\���L9�n8!H�)Pn���ى���)	�?s���1�!^׹#�x��5��k�1�F`�
1�G�e�債	݌b=6�dE1|�wxչ)k��e���!������r�M�xⳆ����_���O��_�!�(i]�x@�Ia 6�E�Q��J��ZG�oIž���<Ӎ9dr~���]�#}�<6}��e�`��W=(J[`�r��9'�k&J�<��^v_wdu����{J���7�RIzTZ��<�(�r�y1��PJ��7.�H�P�dz��!^��C`���SK��K��)Xu��U�əB/u�K����S�9�(�d�7�-������X$t0�zT�����r����B�$h�n?N=������S9�-�^^��57To�ԳeFגh��k�i� ����S�#�`+�/��w|L�y>ˬ�El@ �7��� VD��`TEhb:^�s�)��ۋ���1� �4�&��.�Mƨ��hR�������� �G�Yș���[�b}]��ټ���v�gH�yw
�I���g�Cs�X�.Hkw�͂�	Ӏ�S⚨.��u��4ъ}�^I�����0��ڕ����A}'��!�;/j��;~@UTB�T|��H��
5���niu����֦U�*ϋǽ-�����t�����r�*� �d��c�cn1H|yII�lX��ޣ�s��[*'�h����*>�a"�Z��&J�1��Y��pO;j��}�V�Av�� AH�0��X&]萨����M7q7>ц�iZkp���Y�j�)y���z�o��������K$D�9\#&4�x�o���8���g��9�=�X��gOڡ}��nW��4��S�u���B���b��SnƢ ^�%�!	_�����R�2��=�C˶%�{+��0��fA漡el�~Jz1-��	��n��B�O�V��������ml|��SE<��|�)G�q�4������,�?�P�
�Ƶ6�L!lt3p! 'N�_��Y`�<
k��m���]��o�֣����͘�"�A��'�� $YC�w��0�W�����eS�� $��h*~���r'qjii>�1�мׯ���Ϭ2����)�{���`q6O*���(��A�Vߺ�bP�/E_����򺳴���2nIQ