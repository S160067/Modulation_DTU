��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���,���`�Q �����6�͍	),�6�md|_��n�x�"u������K �5owJh�E��qڑI9����%,%UEwf�x����;.�9��p3��,/�֤����"��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf^��$�i�g�Wɐ�)
�Ql�Y�+6�iѰ�^���d�u�.�Ye�ZG�$*�f�pM��Y���f<���YB�H6]��^�8�G{��:RjeQ��2
�ƣː��5JLO%/.�)����\�
,��YIw_�aJ�/��]b<Q�	��E�������^k	�:u��>̴�_}iT˻����͋ѥz9f��� XnS�{�����#Q���_�=q{���N3!\�w�4ի4��\�ч�����F�ʏ��d8q��� ;&X�`��6��9Sɗ>��)�����Wumg������B�?X{�$�dU�	��`�K������Q�55�+`a}$J�����&�8J��Y���%+V��
��0�W����~k�6H2)L e@�r�1apt�k�������:V���d���\��衷��,n�~�}J�X��atuފ��kLx��h#6��H[�p�B�� ~�a:����VV2�g��u�!H�� n��߬�<rA�坷8�&���&�e!�cc��{��s�G��ʢ�v�]�>�n�yA#ۤ?�F��+����Y]��U*CO�T� �\ ��/�&�%�Μnl�JX��'��� ,Tw�@��$gxaKgU/�k��Wt%��S�v�>#h������k��<�2��aQ��n~P�����og���<�q��^���NegY�W�xv�"����{�5 y�RrlT4c̒��u�X�ݡ���\���ʾ�Vt���bM�ݵ"W�\\�j*�4i�%J9��B�X1�h.�b 6_�k�)Ձ�����O)�����-�n�B�g;�ۊ��)j�Pkk�͎Re½��g,˃��<Iu 9���o3E|��gg���P�:�'%�Ö��c���=(>3�Eŷc]��B����lĒߐ���ۙ���p'/^n��x����n�dTOA��I�<��5à��`L7���r�7sR���STS�m�򕍎`o���#檹��2\\)f��2Z�v�^lOK�1%���-G�U���ϣ����j�_�ѾE���Y�'���V��vȊ����󽰵#J#ǖ#$-{*�/�h���z�t�h�C_��4w�]!v����65�I������_5�tg!�\��\e�~>��~�}s�H��ߙ�s�<��~$��B�N�7��=�w�qZ��#0%c��ĴV��&8=>��q�:�	g6��pw���	:,�}����8p���BjU+W�����0n�v���G�b��'�F*f�.4�4�`T_,�:��P��-�ؑ<,��7�F�t��w�%7w�|�+��'�X@�^��غ��
B�X)㿈�n�^�5��vP�����.�&J�,��ц���*6�u��y)3��#�lm��#�1�<s�7~�Ơ�V�E�h�>8K��Ĥ��6��9;��|�'�5#�C'�݂�I}v�P�u�K�E��8��y�z��&���q����-T�$Ȅ�ޔ�t��P�T~�.`h�Qt]h9�W���f�_�5Ԍ�INT	6�#b��3�|�w����,㞁oG�:�}XBX���"yt�ot'�c��o�Z��C� ����\+��
��[ʤ*,�]pCm��2yn0�_\���o�= ��]�$mNO$�^p��*�	����漑ch.M��q�c ��?-��P4���v�o�1��K>�����W�$���Lq>�����B�C��eߎ�+Q��̪��u��1f;/�2Ԏ(���M���4T���9m`�3n��v��r,US�Ń|�pW������5�Qjy�$O �c��z�ꢩ�p��a��ܰi���2~:�P}�U=�o��3��q���~$׵=��g�҉��q�$���T�. �'�
�D�3a�v2�"
��0Мx6AO�7���P�_�%s{� �*I&�u��'d� Q�;M��xj��))8���QQ�Z�"���	�j���P�����X6 Q)wܻ�%@���a�q��Zq�����6��Ö��S��ɟ��x�W,���ϳ�0�H;����I�>($T�z�<V�ڶ���X�˞ԿP�nH�
��>���N�d]R�c�i����"G�c��\=��~0�<�������" ��9Q�/'�������	�e�F��\B�	�R�Dgt���٪�|E����3[c��A0u�5b�O �MP�8� T�2�zs^A����rn\f�Y-��Q0
�V���O�ç�2Q�u�ej��!EM�ο�� �Q� c�ZU��mJ�=A�b-z�)7hC��
��(O�������s�pm5���M�5��W܋�r-����_)N�|�B���=�(C���FJ%Nb^��̞�5Q.�����0�|7���'1�֐�'f�`����KrCAg�J;F� �:֓l.g��F�X��^*d�
��2gI���[OڵT�,p�O�W�5�V�����͗����E�Ʊ���B~@�0�:��G����������{�6��ӵ�ɫ^�dBa��A'�W�m!��(��q��n�+$9��\]-e���>v�|FRa� l�:}��qz�P,6a����E��E��u ����\�FG�O�����f����Z�	�unWG���i��h��U��V��_|,�0e1S��<��P�*��M�����ݤ)�"y�y��*�H�O�y�9�٬��:0���5c���p�o�95� ��c	�/a �ۚ�Y�l+�\ۚ4h]��5b$L�qߖr_}��V��Jp�=��w���ˀQI6g��Y�lދ5y^�>7��$���d��FO\08<򵩃���Rq��k��)�7���Sv TN0��S�+�[9  %�9� �@���i��fB�:B��R�+ I&��Ba8eB�W�X��F�ú�'��s���)'I�?Sqm�W {j�@��c}Z<����#.�漰7�N�N��we,���y���˪L����7n���#٘`!3��e>�5G�YV�v���A[C��{*����8LM�Q�u5�s�L �Q�������麞;"�e˙�!J��@ӨĻ�ʢ�u��Ԝ�WdUk�-���N���}VB�=�
�<�l|#�����5,���dd0gR{þ����J��PRH���Am���b@� �B�*y��t �I��#������̞l���)wMk����G��{��h7ÞfR�����Ka���g��QWe��XYj(�"�8�+�s���%Ջ�U�.�/�*nB��5f�wo���r^��@��O���p/6"�i��1��k��Sᾒ���w-��RT.�T�N�+�x{)�݄];7�<d���߲�(p��.���NG��qcC}vz��3��l��r����`Sm9[I�ȡ������l���rK��[��R5�g�.M��]^���������ywϥ��hwE�?�%J�#�5����@���0��Z[[mqw���a1>�C��vM�:h�5s����k��^|V���L���f��EA7���2��D�t�4�G����|&�)l+z7�,Ar�p*��!a^�e�ͼ<���O`=
w$t��ɪdu\��P�'�S�I[�K���ѡ�/�p��^n�7ϡ�1D�&W���� ;�H�W�ɖ7m
��Iώ���(��C"t4��B[�����8OvA<�(D�m���Gc�����	�S}C*��w�U�e�J4�����_S�����6}NJf�aQ�t�ᾠ��
\F+�����A:"��2���<�]�]�K�:,�1��d�L�>��ZV7}��M�Qg����W-<�������#�ֲ����Rý_�x5V�s�7ݼ�~��qL�8)�,@g�;h�����}���`��˰�?h�F��=�q��X�/{�޿і�Y&ߩqy-ܶ��Ȩ��tM�s{
�B�vE�(A�>���0b����9��?#������� X%Lh���	"����u<�	'@�h�evs��6��k8����Wĭ�9���O��0�����3MPVSZ�f�އ�fL
������~�%'�~nVf�D��2��bI �BUń���b���>:���[��HL�۞�����s��Ѯ@��`�F��t��#�!k�"J<�_+Y�qG�*���.��*X283�6����]A8����VA.�G;��:�=!�ķ��MB�S�NJ�3
��>�?��������@
�tvƱ�����~H&5*a]�`�:M�R��)Qg�i7aK(���4��Y	���p�����Ŏ��d�g���\���6r��;��\yW}	+��3�7k�
f�ǽ&*��c^�C�ѵ�k�藎UnP-��i������`����U=���V�k7A.��e�7�	��z��^��9G��	n��ަ�d���dQLRg]>`��;�5�#�YN)Mf�L�6ɴ�������ɜ�H"�1���VZ�x ��HZ�#
�~)��v����+O|���Nh��g�#�S��7|_ê�+�֡�X��MmB�����R�z2�S��Kb���|j����v�tn�3)�=�y3����Ӈ���*��H�%]v�F�� &hԜUF�6��̫5�:�j��	1fFc�2��K)�I�g�_]+;5fEx,*������`��ى�3�Q	I׉�5툡��C�IIs�w,x��������bD��+㮼����x쳸����Q$K�L����\f�O?��u�\�s�����"m��������tN�̔�Ļ��q�ϛ�o����w�#v���$��S�X�9���Z���EC��~�1���|��XNIMXl|r�U����:�g��g4W����b'o��d-�bw^Ӏ�!�Ye#��H Fuc�5��p<4Z�ą��Ki���$JY=p�~ȗb�/�-��	��a���Ĵ�B?���L+�|d���%����%��D`F�̆��6�@�Y��t���̧�]턨�Qmu�um�j/�����t����H�I-�(��LH5?��,�-2�'��.�$l�,7sه��s2�g�|B�p&�Վƛ? �����M�����i��`i�8Z�}��>^��h���o0�>B�1�5��NצlXYPc,=ى���T�Q/S�r��F���Z!k��<qL�|Z�C'���$�%x$0�騶Aq��O7�f:����_�=�b�*��]�c����-g��*��$`α&|]�r�0�;K��qſ�I�@}��χ(o�*G�U�>�:׻Ņ�K�u�9L�F�X �Uk.���#]5�ZH��ε�3�g˯����f�$�G�w�摧�"α�JO���B�?^�qa��7(���l�d�ty9�g�3��C�����<J4c[�kya�f 	W��("0��z�F�3�)���9�.���2��lI>�VY��to��������Jc#(�R^��;�p:o��&�9��w��P������� �F���-�1�Na����2S�ϩE������8�:,6	�<���JD��+g��F�'�c��At	[�"u]�&Y=��cŧ ��o�R:ǩ� �8X����2� <7&8��0/�Ҥ�F3�����:�k�Æ����)9g��L^�N�'�S�?�[�v��Cq�	y�|=y�ȉ
� `Y�a]�康X0Ӌj���:�"��%�VYQh��Q`L�>��ٖh$:R(��	���56�`�a�t
OHaܶ�y�#-i�zP�7[n�V��q�Ѹ�%�4�B�I߯�lH���DY^+��s+>側f2��M#%���� ���K�7�!u�{}:��0Fuz���3�kz��Vĥ@����/��l����Y�ń�q@^K���5�ƥRuؼ{����J(-h�W���U@����/��Xΐ S���|�wC�c�\R�0� �S^��d�����	��7����Vo9Л��4�K*V��N�����V�,��XG�pKx�i�d�=��>ȣ
R�CHj������YŅ���ژ����t�Geh
ITfi�1�`y����d�c�sw��1c��4��k	1S=�,t��aq�[�E�!{;�N+�֞��h�S�5*'�	��D+-�B^|=�~nZb	+FVGM~�+�+�����?iW4�+�E�0�U��MHC@+3:��2���Niy��)��vχ��t�x���?((�z|������E�:M=��Awtv(���^-�R�"艞I�">�^����F���
�P�*��n��I3	�x�)����{	ԽwN�{���(�/ʛ�����O�ý�)}���vaJ/��o�ɱ�@�H�wM�Ϸ^Xw�����n��]&���i��t�b~0����HѰ9D����My�1+���k3����M��Q/d���h��r���r�� � ����\��Ev,�7(:}RT`G<"jQA�+��Ka�2��\O��$��k�`x��6�D��8��;W��׸�yϜ"����]��{b0��V�G��|�[��
�1xw��)�!LU��Ѻ!�A���K.R�fj��8�T��騈rʈ�3� �.A��x�uf$��M��aQ|��{Te~Ϡ�����@b�������j	�` ��CR~F���C�y\�rDQ�._������Mk䨌<+��������� )Ȣ��$U������[#����Hs�j���Q�k�i&������7 �rʔ�T⁼gE �'1�����3#�L��^j�L��ju=���:&��mR�	�^�s1|:ɧ�yݹ�����jC����{���G�OyO�OZ�υ���5�Hӳ|M�.�ez�H�|�#��_Ż#v{�\uj��@�m�%& of͇�eKY�$\�''�/&�z�3�߀��w������G���j��w�i�L�R��[N�Ȳ bv�w�m3ZHw�7�P�ȏPUp�$K���:cN���W�ꩦ@�9k#�(<&P)|��}�\����̿U�㼃�Q��yeݮ��ٛ����ab�m��I?�c�����&�+�Օ��O�����51;�li���9�b��c��&��pl1���w�����B���g!�r��p�U��޲gy姧�L�5mL@�]���!�j���x��uKl��&+����'Z}5Fq<d�28YW�w&��Q�'>�7�'�2�)<[E)Be+X]{X��~čH	��!�EQ�������CE��)@��"/ p��|�
���wq-��^zoN�T|�!j)Ϸ�2�%�߮J���ӭeG�x�~yd���S@�Y[��J�hr�Ʒ��/�ŪJ�K����C��� ]u���"���xƴ�v�$�߸_�ˮgTʸ��G���	KfaC0Z�|W��� ��$��Z�U��s���8pa�(�H!�_�}m�d����_�a��`/�ؑ�{�!$��1����*JA�l��7�Bu�*Y>wK ��ih%�Ŗ�x���m�Efw�(#�\���ס������U�4�|Ƨ>?��$5�_m�bf����N��QZ�t�$X�['ۍ�.�pC}����f5$� $U��O�*,F�:w�D*��ˡTig��qm��T���a��7;^K����V�6�A}�u{S���5hĽ'Tc��g��N����`�ȡ;q��T�c�ɱ�mh'8�#�Ks��BF��}&hC�8�����\��"Q!!&� p��oȹoҺTc��܋D�T{�7��6��i�l ڶ�}�s0&���ۯ�qky(|Ν!�l9�G�I[�Zɽ3�)'�;����s$_��w���p{�n$��'����8P��Q�m�Q�H�d6�Ǟr
E}Z�8*��c����kO�]����g�,]?E��;�����^�)�=N{��j�!�':	z�R�X�x�Q�	��E��=����ge61t�t����S�����5�LXp���DYZb'�0p �+���b�ND��bI�T������Ҕ+����,_�1#�t�|�.bZ.A{c�2bGV�jV�j��w5�c�KV-��ۏ��TG���!�c��^��(Z#��F�I ���Y�����'����*�rf&)�:[�ٯ�Z���B;��r���E�����Ug�$Y��K�3,��Wһh�:cǢ�A�^L@$�������(g�*�R��]���ąx�˿�c �<�sJ�g�_2\�3�^{����Kr�z���m�:`��5��Y$ʬ���-|ԏ:h�l������V�"�!����m�צ�]�PGE;>��,|����lx9��)�OnǶu�!K�;�l���G�~�����go?���鼕M �gL�w��abo+�c5au����](�S6�K��t����k��-�pa`��a���1���f�#�m���E�l���eM��tTX��YD������E�h��da�v���O��ͤHYz�uv�68k��Y�6�����)ٛ/�.�G�w�-N|��3��1U.�u����C��
�h��SJ}�Į@����9��4���xmt�m3{��M������7���+�;��c��ʷQ�9�Q�C34�+��+'2���Yeު�=��#�W��+{��;ƨ���Y!c���sߵ���IZb^�S���N�՛��	�^�Ѕj�s呗�=RI����#�,�K��G₿Z5�@VR� Ȗ�t�8-���u�+`��Ϯ	[����x�x���Nv� kF�����6;S6	�n�,��*��&��y3��kdde��Z=-.��WL6~m$��W�2�S�_�s?	��"��$?�;�����kD���|G���6�@B�__�f,�?�ץ�׺=�����1�s�pwTj�fz��{������M�O󒈕�u��IS�h�ɮ_�_0�� �A&�	�^����1zQe���-��.�b��􆁽 �;����v��8�dǈ�+�*�����ĦV�8=;V�3�퍵{��4���[���H�l�wي��}/���y��L�a�GY���\��jz���^@ JM>?zdJ����������S��h����3xr_�l�و7���W{Q�I��wk�XJ�bR���Xl��r���#��d���c;��M���8�wz&�T�+p��Xh]졸�e�������V�bUxQ�����Ez�x�WX���8r�4����'n�9:�U(m�^!�L�?����=2@I���7~�5>z���ho��|f���4,���{;��>$}��Ͱ~��Ht�L��~�>����x�GS"�-T�hr���~�е{�StNSZ�6u^o�tϞ��͆}�B.,��� ]I�Yd�f³�(bH������Y�,��p�
��,W9��:�v�=%~Kz��:f�K|ǘD��7��uV�x�Ɖw�է�kO�Yυ-3�x/���F�Ϸ�O͗Ҽ�����0`  �X���>��)���~�e}��\�D��m,p��?5�;��JNq�8�k�ɧ7DV+A*����oi�]g��[Jb���e���6c�Qp����sFؾ��	��Y��;KD�NiR�/����N���7��!�}�2�};��N���˗*sc��n�֩�|U(��iA�:S��C�¼1s���Zy����2����k���5K'uz;����G�}�}@�Y= +9��[n�������s���˂0���5]ݫAX߉�����%,p�fO�"4��TMgK|"�S�~�y�]����\�kR��$R�)��<�QCG�4ͦpK�6�X7�+u�:5�ƃ3�z���v��֩�岂D���C>�w��?��XY�-����bw��fԉMo�{J ��Sf*�J4)jBE7\l<�C�R�=����P@��5N��]jQ^2B��S�70/F���V2-,���e|1�9l�$-WM��l�ᓲ�lj�R�bSЁ
����ra��ܸ��aIM���S|P�S���\谜�������4�:���}I�����!����o���� J������� ѵ���@�}�̻!y�s�Y��,q����+\|���E����L5I��?�D5�p��4�!/[v4s4�	����K|��g��I��'$?-�W�j�F�2�VߊJ��r߲M(s��v,��\г��ʤ��-������pv��Mu/_��H.�<�f�CC/��+ßUN0����{��6U���<p40�U���}���lۊ8ּ?��k���^pv���Nv^6�n��Ae%�j|��Bv{�Ri���OKJ�gJy���4%���1RǠ�����%��5�d��
�I3����x�Dը��%3 1m��S(��>P��}�o ����I~x���f>ڝ'��`J$ƨ�S����i"
�x�/��`-[��6���v�Y�:l�f�[!�4g�n���_�v�)X�8m��Pe�3}(p���JC���7n^��6EʍhR�m�QG).@�q�%�ݻ!�J�Ӽ���ƪ7F����,�*�D��{���`�mC��	>a���D@�njyJ�gi�b�ϗL��,�j�ms�M^��`_�D��z��a�0�e�;�l�n�w��U�umU�@��t�](���<��#��E[�6kX��u�Յ� h��f�9C;�#�3T���m�1�d��O��y��R ���Mn ���-��F-��0�LRVT�4,XO��6�SpW�13�=)��sG}��D���͉�ϖ��D��Lޭ?�Y`!��G��g'uY��z��H�E�m�`Ǯ�yا�X��֝*[�q�������4_mt�ƿS��r�-�hGHwe�� Ze�
aۙ��x��I�5Ӹ��s�0����+�]�2�e�?u@K�p�F�50��)�aZb���`�����>��o8'�B��3'��8N��e[V}���>�q��B���f���������\H�qN|]���j"MY]��M
&��Jf�1P�<��ì� ��_xW��v\��ٰ�wBN�-�z_��z�l�;�|�a�@�?�<����ˡ����\l�X�1�+Mp@���a�� P�hz$���$�2uP�z
�i��O1�*��{
�t��RM��9�/��/R���"*D��{3���F���K��]��M�	,zK�����"�:n�ꌒ�.}�wH�Ǔ�+���j@HW,
����/��NOs���$�s�f`�/���/��c
+��e�aMm�R$�1��S�[�FAx���S���ѺI��0����y�z������e�HU�S>�K��b�~����Ld�ٔ����@�����T�7�6��e �#h��48M'%=���oE|MS�1]����V҉�����"��&��Vϱq;1�5�s�{�ۉ���swe]7�؅�b��G�d,ԣ����S*�"���!\W��3f�����j؂zv�R����YF{+4{XڥI�ٛp׊�=͑u%���7j����|��6fg
[���������%�W������݃�a��e�%�g��/_0\��ϙCMM��J	e�%/^�Z-����V���^�b�p�)̛�^�yw��-���j�?����rˀ_/QN��1�����x�p�L_X�!��\S
�c�̮�n"x�R���� P�2s���aK��d�L����� ��Hu�m�w��|�=��0�)	&	���LMd�Y�`2���p(�� ��`��IMljN6lH������:�AH�~�	�p=��K�cH�Nt&� ���m��x�G��5��Ix]��.f����o8S0��S0�yEx����5�䀽?�=�R�f��3�M��۪|����^�.��'��J�v~i��.��X�q}�l�k���%3��0.�NeR����D�z�ji�� ϋVk�����
b�~tU�q3���c��[Q�J*��.����a�i� gDp�F�&��	�����׮�-��8����ދ��D�o\��0I{N���"?ß?�͂|Ҧ:S�,p6^�r�I���[00���p�Q����]� ����{���K�S_	���(�-΢Rť��/����{\b���
�2�^.ĳ+&���\ϯgY8#�y�\Om���?�{�D��+w�=��ĩ�,�y�)'���XL�b��9k�U*R|ЋI�����F'l�B��S���� �e�``�-����#�$�����P�%{����8D��f]R�0�z~�"Qg>FȔ ^0o��n'�;~��� �n��H��U�)%��������^\t�qɂ��T$ޱK7�BQ66�	R_�]�M�q���Z�����G l_��XL�a�0��&���@��g0����d�->����C`#����0`�s�gO��� :([:��z���F�0�a�z�>�Cֶ�Y��g��p@D�8A l`��z3.�Gĝ�g�p}��y�<�qOR-dH� R�,�����ͥ�Hw��:���Q7ݘt�}C��Y�����㌂l�,��vA�Gw��Η��R����m!2w�2a��X��@�ףA�@��_�ަnb�a�Sќ����O�S�ν����@J>�>k��nJ����KGL�X��Wqn'fV��s��ۂ���$��Ү�rg��mp�>)�:X�]���&}�cyFS'Ѕ�J�30x�G��ZP�ݎ��\Z�����CT�G�ХƃA�L$�9��~����7��o�k�((=�b�W�-lt�T����D��L�i��X��IsT��E�1��@3�ذH�,��/����ޒtJQѳ|���<�כ�"���KW��-�3�cg����^)늧&]�f)�z
o���Z���Ps�e�BТm8��k���hI��1��,1@4!s�Eݔ;�"p��H�>1�J�|Y��!��/��W� ��7�����F1�}�S�����g]��(	X��!u\�1���b$/4�n87C���ר�5$p���d&re���WT�4���դ:�MŶ���D �q��A��~��Lx��!�JCLue���I�#[�V���M�kz-e���bS$?M�&>��N�x�I�(&������]�˛�S3C
�i28\��OU��e�x����Y���Wx+B������;o�z���(q;!����
pU�,iKh
S��lP�T��4b�o�^Y�ڧ��3���?�A:�?*��Dn/�?j'�� �(���|�:���5�{�lޤJ0�HO��c힫"����ZB/|���u1εv��	��;(�ǫ�t=y�D�t�߶1&ۧ/3�u�������yW��A(༏@-��|�˿�GGxe� ��_W��cC��'�eπM8�̎K�����4x�"���\��:t�[�cm�گgJ^=��*��Pb�邖�F��n#�*z|�3�R*�҉+�ЇX�OÜ3��%��5u:���}ER��g��4;{���,x-/�>�u�������2�b
�{�^6��q�ð�� #ao�g$�2J�8	Y�[K]a�g,�\f�A��oXo�DXHN^��Վ1�?�R$)F�>9���(�H��u�� ��1UC�73�{���ojp���p�w^>@�0.�U1��+.�@��8�^�.饧ʚ���[F�gXܿ"��;�l�h�Ѱ���� suU�m�y󲎈�Vh���E�d���2���/C[kK�R䃗S#���\�Ĩ)j�k�}F�1����3�<7US$3lKX'4lO�r���o;<�DXlf�`t6�T�d����k��r!5f�(�l�צ9D��J\���^R�
�K��`�h�x���"��9,����u�҃�J��M������<�
��P�>�����%c#��hj}W���fVʊ�8����
s:�G �㝬�q���.P@81���%-�Ä/��^��(�f;��u��0��N����*X*-E�*�'c$�7y�!��D�Va$�ʩ�\?�lC�q[��c���ʛ��=�����ɯ��"�^:��ݗ�z����Ѫ�⽎H^�ʯ��7������N��D����O�S"F�؟樇G��|�w�u�&����>��^)�U���~�@@�A���M��gM���[�( �Ѽ3�����>svF.���ƍ*A�H�°��		���
/`�N�o��9G<C���_P�<^L5p�]HI�~*^C�����!�(e�8�1pF\{G�jaѷ�;i�AU����D8�9.va,c��Q$��_���E�KXLIEQC���p���z:��y��'s��9�"����;2ڍM$Mj��lQU:V�_��7�Z�(��H;
���`�Kl�X^�n��8;�;�P6?6��6h��|Ɔ	�m&'�@�U���ۉ����`��4���=���y����C��x֮�M(Y���n�?�1]��I}p�[��h�!�/�s�ZJ��D�W�{Q����%H�P8�`�6,aN�
_���*5�� >@����%W��?ߟW����_V�����S3���݁A*Q'�0�4IW��C�d)�8gm�Y!f{e�-,, ���^�n��Z-M��{�@d�������eۭ@��JQf���n&U�.']uX��m6��xo��Cx�"4=�J��Ԫ���C�  �^���W��ãcٶ���B�j�6��ا�jy^5 �E�A�D�
I}�a����4��o1�-�@�����S`$�2?=�m���b�l7B�M���N��f��N�Թ������T�Sx�m��;JsA^�b����2f0�e�+� �G��l)��/�<�I���z�zd��f�X����
(oD��$4g��TQ�)��g�ْ�E;Cw��Y�h=�� z�Y��n��+�T�r����?�'&I;@����{����U���c�3�΋)��F��6�S��3mƺ!o=q�#o0>���-[�l^�ǗA�Ke�C�:}L!4�i@6�+�g-�G$;�m��*�-��G�xC�곛X���&Y`sl��_I� �������u(�喪���EJ�*���7T�v'NJ�9d�n�7KT�9��9N�q�h֗��Zo���?G�/+��y��b�;y��=�GH�{s�V��Jb�>ƥ!\zIfk��=D80���n�7���O�������T;Ȣ�o�T�ܐ�Ct���28DS��]4��z�{�[Qf��w���~�a0�ggE6��f&�4�Y��*+�j3JG�S�u������
?��E�EoU@�_B.�B/$�����Y
�.��I,:"_���*��;�C̹i�"���M~J�S�Ј�|�<�5�;a�!啰V	d���l�o�⢕�r&+�[}Z��r��K��y����F�C��-�p�_��3%�=\`�]�������e����9�s|*c�Lyf�Y�D�I{�t=h�},ǋ�R�s���ħ�N1�O�s��(R#����kZO��O��X�������#��p0�qjh�K�A����%������tE�h螊�`��ܥ�4_1A�NE3<�FW>e����S�!:��O���-������j��@D�^]���$.V:7�0>p��6UK�+2/;rwZ8�:yK>a��[Y��)K,�Wa�Sm���&��ZE��l@rb@��ZS��;j����� u�5���8� ���N�*/��ڴ��p��qrs�����ʮ%��"�_���y��}E#N��,�NoS֜��{\�aZ��Oq�2��K�y��¤���!o�ze�{?!B�)�.���J�?]���Knli�# ��[�~E�n�{PJ��������,Ӡ�	p[�NE�d���?���A�$/6�+��i
%�3��C���N���S�9�IV���#l�̄o���Z'��a1V�3�;-F�F����?������r"�a�.��A�D��C��/f9���9�iCi<&�ϫC{S���&E�\����B5��n�م��Z�WvcK�I�8FU������������a!�|�,�����%� ث�f,Z�S���a÷��Q
���k
N'<�H�|-���w���MvӦH��:���S%�#�T���{������v5%?���O��@�ۙu���KN�:��u�s���C�x�KXB���$��$����n��D�i��i�?p�Dj0ι���W�xF^o��B��q�U�u9�l��.U�ʓ^ ��5�`��Bi���I��:R�fc�dQt��_��?��p3���A6��3�-*E��e*4�7*s��Ln��/�#6#��t;�s�UP�:�y��&|*m�m�r�Q��4OyB����Yn`R�@SJc�{���8��Z"��I���w�2=\���V��A~���K��c8ອ���c�Ae��ލM�;5�Q��w�h��w��fГ��̥T�m����}nktهQu�K��_Q
@��"�qhD��q����y�R�Y�[�!��t���u����W%pB����G�'D��Pa�/��>�ЏT�^Y8��MA��º	M�?g6;�?�3�-a=½W��"f4xM&��f�%P�s�:\f��Y����'V��i2��g,���&d��w  ԓ�JĹ�t�@���b�i<*C��m�Aj�0��L1v�皠�c1YEn���� ����6�����'���8l�ȋ��WS�B�b���W���w���hi�b�t魖pYړ9�[AI gJ�$��ED�egVN7�D�5�v	[����܀�n�@U���6�Y� |TL�5Q��d{-�[$i�v7.$���dԶ�8)�v}Tv  8�/=��uq��x�����2��������xHb����ᖿ��@�{j��ݠ��R�J	s�X��-G<�Ccӂ$m�R����1}v|�i?��V���9�ۯ�:�������[4w1p��V�:FU��dDA�%!�!@�":$�SBY5��\7�S� ���n���æ���®��$4�E-�t�S+��d,Gf+pwN�BP1����O��v�IA��kC�r&5��Z�?b_�[J�^(���\��7|3,Ì=�Y���=��x�����_�Nz�*K$|i�$��S���8�F��W@Yv�b��*�'Ĕ��>��>�띎��Y��0
J��DH}e,��1�N�f�����J�� ��aW�'��0Cg,���[c�}W ��R�o��-��a0av�)�J�*��![F�x��ԇ��|�xO�-M<򐍅z�#{mf��B�>�}$rK��V"Sv��Vl�m�o?>Փ�Q[Ɠ"TvI=m�S,��J�!~�&�mX�lo�=��$�H��wF9jC��#��:cD�Eu�����v�K���������qY��u9I�ה���C��%0Q�0�'N7|v���ez�84Z אgb�U�
�kjS6���m��W�Ꚍ�t�"�t���,Q� �i��h��� �t�h��3���ӑ�Q@�N�⼰Q���e\��| �������#g�'�3:W��=#B�6�lb�L�n;3�]b�����ꔛW*=��0ňJ�Ti�>Ӂ�?w�.�a!S�UZÂ��l5��\ H�����ZO7����Yf�Ӗ���\��_�E��2�Ld��-��!5|Y�>��9@���Kc�7���d�
w/I�i�>"}��`�k�^*�9������q��^�7��e�o���Q��X�p�m�v=p*~},�����3�^��: �U���y;����G�=L�t����yT�-Y=*����QLAɡ�"*��B�*�m� Y�����.r(��W��Y
�=Dq=�)�v3�&������u�����͠��򃤑0+*	���aa-��r�8�8�4O�cl�I=�K��[c���T
NZ�j�"��T:ѰF\[u�cP\3m�5� :y�q��
�E�#��nyT��l(�3+��@���$�F$~��Q
�_�,nMN
{/���% �ȍ>]�RH=�R2���
?�*���S��z?�v��C�CWN�[9��懖���}��7	�Mp��^S,�4����
*|m�䎄��Ƚ!k��q�;$8Ͽ�����d��Uv���8{����s@�?�~,W}<1�vHlk)�@����{~2��4,)��F@��vfVV�ɘL�B�t�s�t�+�6�h~��87����T�ܖ�#��[��f�SO����'fvg(�=n�-�R�J��k���YY�W���Y \ء�=�1��]=��� 5:��Ӓ���-�!	��Ů�%�\S����F��L?�fv��qg���Y.6�:-���}	� ܫ}^�A�+��k��rv��$M^U�$�#���Q�D٧�*�0���3(���2��rqcPv9��x��kԊG�^(�	�z&�`Z"�4��b���LGO+�)^�Gk���T��b:k�����,o�3��rpL�ϩ@����Z��FI'򻸫��	���n�`|�H���� Zr1��'�@}T���6� ��W�jJ��DT�-7���X�rǘm�Ú]���ƺ
���^��k�&�}��*ȇa'H޲ -��8=+49Q��t=e���3g�a��T��fY���g�B�Yh^)����A�]aۓ�������t,��}[�S^�����U�0ǣ}���j �?)�요��QГ��.#ږ+�௞����q��C��5wW��M����Zsz�&M�'�5�:̥�̆�+�z�_� b���,ᕁ��a��"��AJR !,r��̟w�*n�0?�1bf�wOy>^~�]���́��*n~�gO}���ׇ�D�!i;�3.azo�-0%^k��ݕgm6�6�O����}��P�G��H��D<�8���M/1�:�*j�zWtk}� �v,�:$��Ү���7�JShf���h3�֚�hS3�<
_�~?T��q�aϩ�­���3�҈3\E���� '��^!���e�=�H��+R- ����8��Im�����]-����Z�5��ST|^���4�J�a����:��2ӿ���Y0�LB�r�u*AqN��ۀ��E�"z(���ct�Z{9CA�XX�%�k�LQ�/�J��=�sM���p����?����$�й���I�c�Q�ŚyBt�
��A�	?�R莝��#�;�7e5�=���<�ju����=dY��l��@>!/廎���ڹ�0������n��gtYP׷ZV�`�T��G����W�?����|�wX�A ax|\���
v޻%@���ݦ�̑���/�Kk0���~@F���屁�;�7/uhC�ܛ����Q���7W�^CS�FHNZ$En�SI|��"�5(O��| ��=��]�fp��e��D'�a]�PSfw��*k���",p�X����,�����L��n�z�>�w�r"�X��b�o'MD��q����+5�	S�M�H
0�hU��$�i���{^�KY�.��;�$�Ls��Lv�P͢�Qx�T[�2�����	ɲE�!i�û���A��I<~���]�j�z�NGK��gԭ����Z�8�O�$���Z�ѕc��p�j���� 9���h������H*�ˬg�#���d�6���)�ƂJ/m����Q�I$�DYs�QwR�2i��*�PW��/tpӃH������ܺs��6^���{޹xH��*�̐%�k���z�����9����	h������jb��W��.��0S�߫^=�t��+�ۿT��B⫗)d�\��+5�r�w"��iY���W��}o��['Z�\Ӎ�����kv�L}/?��wN���0�s�g������&}��j�xXd��m�^��7(�_w���?����з����d����7>���	r���b[�/�y)��Ӵo{�T�ecA$�F�=�Ў��d!$& �e����k�&@o��ߞ�ƺ�R^Ǜakߠ=$�>F��4�<8ԧ�$�$Ɉ��x�e���&������p�����K�����I��H�U���-�C�K��M�,�l����P����73�_�n,d��/�h;���9��&���ؗ  .X�ޭ���
5}�ˤ�U���υ�w�txmS��<�
�_��	��%�Y� =T��'�ʍ;���r���%��ţ"������{�SD��I0�6�y�c��(� jBS�:�8��s�?;�(��d8�VЖ��w=����=,��WBӤ�n}�1���j���X��t�����Ss��jǮۼ�3�),=��K��;Y&T�T�7�K�+�!�+�3f���͔׿+��j�Dq�yNr	��F�Ǣ>ދ����j-"�֝ϼV�����KC"�9bW�%���TC�:�z�5�'j�h���
[(
�tڟA_�CC�^	������������26S�O��������<�h!�FA���SO�9�M�#�)�Q��TxF���_E���vЗQS�뼣,|���%�!T�]<o�]>lv�����D�\�nY8j�@�����4�p\�A��<�������&��(�}���@���fT�7" 8F�P���:�n6�!�'(�C.���R�Ǘ)�E5o?�Fxsd�_=����Ш�9���^���)����8O;���M�Ƕ���9��5�O��{B��;��!)��Sl#zb5nV�
�]	�;'1����K�'�5����V�I���\�\V�t���!��S;:�����'p���5}F�+��,�RIӹ�J�� �ᄣ6�5r\���2�h�2jV�4�Bb�UP.�L�nD~��L�3�.�ˏ(�Rֿ.�]Rbg��@��u�v��qL)�\P���8��ڍ*y�����9�F=���(��З�چ34��,�sX�X�ƙ�ޘ?��������q�+��}ѱ��l���Q�
!�w)��~��@��!aKa~�R�}I�~y�e�R��!��
l"�w��^>!MgPρ8���Cy扁����JQM����2�k����P*+��e���CS^諏�C�<��O�rX:�b.~��wA��F
8��ԓ�s9*>���@��"
���36��%�>~��#D�ˌ��bmx�$VӯT��]������p�p�\v�\�2ܥUH����W���d���	��UI#�ݑҪZ-Y��%� >�X�F�ģ�k��������a�Ù�"�";�lxY��4C9���!�e(������h�
'H��\��W��>��O�Tь�J��c�%[$���FѮf�r;»��^�F�'���QwܟR���	��+A�Q�]_��.�&��#H>D��#��jl�k����QS��<��GEJ{��+�j�8ԫ�������ʄ�ݮ��&�z(�t�Rc��0�����J�o�ٰ�������b��	0}�S���m<�а/q�(t1Ƌu#g�j�pC���4޷�n7N�f��LsS��S)�,��}�2�beC=b�/�ț��b��`$��oO������B1HJ+O0���u���k�1%�ͱ��>K&h&��:�o��))��:���֛B=��o���ej"k�Y�2�L�����q�I���J)XO\U�JW�LsvmqKW���	��j���P��r�VN��d�D�ƀ]7�9n�?�iw�"��.d�BR|��|���=�к����cJ�R��ࡔ�~�:�teJ�մhۋ=u#�gz�I`�r���ٷ�95�,*'�?y�.��h|�� ���9��#�:��h@�^��5��
�o�J��
�����Q�b�:��놗�Fc��8'���TZ� ^1K��[e�5�֌`�!��A�˿-����sëA�^�?ƛ'=�PɆ�|H�J8U�77��W���A�c��U�胙��P��wz������.�5լ���߰z{�8�I�ә~|+ŘT�(�?ۚ�Z���-�,�ؘJ�X�(Ƅ�l�s�����2�ŭ��k��E_G����-�a��L�:<�=��4'z�t��/+[��.*{D#�vF)���ȼra�R �Vğ7���g%�&��)�~�������?��8�}� "�&����f3�%�|���>��SYc�]hסj�/�V����Q�EF�N�㣃#��/c�.9����;��Ȧ$7�SJ1!X��87�4,|���'j�%��h�N(�_�	�*
9�L��oz[G]D��Qh�v6���|@c=b��Y�0�ػۤ����Y�\���C�������=�:ʳ`9���+�Ѵ�o��ڛ�`��j5uB���<�,��|�l��Vu4_ug�\oP�0s�7VO��B�y5��ҍm�~��uF�q�i���\h����-|�B��K����������G����s�GQ_�� �"!GH��u?~a�8���TSo��u������c.D5���*�N�>_��A<1.�]��7��ĬZ�$QWb6~9�he�Á��`[)+=t�W�K�8+[V����?����e܈��r8!���4�� ��V�SJ,���T�\�C)�.�o s�^�M�1�O���1m�Hw@��dI�ik�L�H�
��Ħ���M�3Ny�T��%w�Rb�;f0�BQ��+Tx�V�\��Й=	�	��Ŝ���t��b@-p4��K��9�7�P��*Q(��nH+�\���Z������I]�H(,O��b'ؘ�	�L�N��H�J�4?R��y#u�PS����*�t`��  t�NLu9�^Y����5;�Z?hb�������"���':�[�7��^�fwϛ��7��}��g�8�U���ͼ�o�C *��˭���d'1$1I��6��kpt�j��K����' �1ˆ���+A:Y�ʅbD�E'<�)�ǹD�H�RnC�c�uo{���d�5$}i�9���3ԅ7�ǩ��7 J��[��ژKV��*S��*=L2H������8��5�?@@���	G�  �X�v\��� |�{���F�k����ӝ5wl�-�'BR�53��&Y[���?p"{�[t�d��Ȣ��@[�P�dW��$��wJ��+)��H � RK�e̖��dd�g"P6Ȳ����j!%�P �nhiI�����s���v4���/�pu|x��f��F����F��mE��7�G[�(��Jf���R�NF	I��E��� ~�N4�4�e�GѷpNEi!����Rx�u"@�0�go�Q��R*���ho͙����_!'� �x��2����z e�v�|��>���0Ӳ����ʁ׹��_I�$�b*bF@�� �@\��U"8����yg�CTy$I��_�<����-�L���k��L�y�99�'���O�d�klft��/��g+w ����z^aE	��\�V�dP� "Pj����@u:{h�ޒ��<k6������m��l;a>l�6��ĹiI�f��T�鰙y����o�I��C�z8TV#2�Q�>�L�C9��Deo�0�U�C�,7�5�o�X	�S^�U?��ZF+��W�����5�iD�aR;,6�����]�{��b���2�a�{��$*W���H�MY:�>*�	]-'�\e��-��o�H&h�nK\����X<����c�b�0M0��!���Ǵ��@�����k���ҚL��i�D�B݇�ʹX+y3����3�ż=��'��d��%6ɛ���?��_Qڊ�S�о��b`�f�d���h��������H�sik����!�-Sh��t(b�����"ҟn��� @@$��l��gJy�����]D�Z$H����1�`�w���`Lx��������B�e��dF^	��4����K8��=F��θD{�@pibH��:Z��oA��mA� c�N����?�x!	��S~�
��A7q��'-��~Y�LV��xU<9��A�`B�O���Hݾp�5��WWQپ�Â�'a9M@@XҬ�qE-�4��5����.�\F�T�.DG�����Q�f|�Y3�k������8�=����,��ێly6r����sNp�� �����F@6��Dn�(Q�L�}&p:��P�*�{á�H��Y��\�G{%8떍1����� y=p�+N1m�$$�N8O�r7A'���+��@6���8�˯ܫ2'�� ��"�#7�J~b�4����y�:�tBM�Rw5�A�O���&����QɫN|`t$�gY����I
t��P��f��Y�� �ݦ�$ɍ��0��~������*�<?U�,�����B�d犏�vf���$i�埻>YUB�X���6��۔Xg�w�\�`f�����k��i��9O�Vy	q�~����ŧo�@%�ғ�㣑��+�¥Z����
��v��F@�.�(,js����R��֘�Eo�,B��cAF��Ԗ.�B"宓V���E��]���س,�"��m^����d�i����Q� ���iH�FM��Y-t�6?�x�)��{��I�9��9�݋���Y+�Аa��Ď�ug���u�߽�lłW�uq?� g�\+�?*�������i�gAt��K\6���vUo6�\1F٣W���0�vU^D���m����#=1Μ^��aUZ8���C����Հ��*��5���G���:'�?5�������>���X��fY�{g*(���ű���o�v7�?�m����N�~�_\$+��Jҗ��7	n���o�0p\[��]�}�f�)\ò�!�0~#���@@�#�=����~���Ou۸��GPb��t=̞���͔��`
W�dC��O��bM�����DO�2!u���M_���U$.� �N�/s�y��F�|��1��co!��fX�xc��gE8|?�Qv��(n7��=����`U�N��_'i#�%f�W�pj�M �ٓ������ȅ�{f�;L�=�V�|�>(|Y3�]�Mݳ�5�d�#��a${�X��FǇ���	�ⲏtiW�J���Pi�E�G�-��F���
�SKJ����K�#���QX��ޔ��r!��vt��d�i���u�}�*��=�-��?�5�vFx{N"��>����o�W*##����C��p:�����!���~�2�wgB�I���D���;����j �k��Ў*;�`���2Ϊ�J�Lx��p�v���f�B����C�Ӹ�@�F��M�ufȹB�|��u���a�ִ���b8{*&�P��*rH4���	7sO�gE�����ٛ�\���N�]��qm"��l������J]i =-�J�u��j+F�>��^Œ��~�#����4�Q��A��%=�7�3dS���Ф��r2�_��էWQ��C���>t_���3,^(B�:�[P�cŭR}��o�ɃE���-�5V�Ox�Í)����h{�Rp	̔�4�N��.fB�)ֺh����'o��$^�S���o,ؠ���`�h���,��*��ֶ=,��@�Ӷz���u1��[>gw��� A�tl��ˍ���"3��X��B2����] #qc
��Ԃ~����`8��D�Ä�,jZ��� d��8�jv����垼�yJf7L���+x)e<!�	7���HG��V����#����}8����ܴ�|��<�H�ܺ��i�d��鼆K�>�cr{#n��^���a]n�p_y������)a���� /�q���ah�W��+��QV�iH�yU�ء�S']o�x�M�s}'�G�59'������<�-"38���塹)�V�E�+'��c)�WԲ�=U��!.�!+L3���R��I�� G(nq���'���ص.�@�o����.�� UDCd㤻�� 3z��S�h>��ٽ+��	�˔�J��Zt�xfqΌ�x[�@���68��H�R�w�N��lMaQ��_>����]-�Q�A��EE+�	�r��5��<ɋq�ԂcdB`������V��#uixw�	��7���䷸�36���b	�8����X��tF�C��S�oX�|݆9�'�
Yh�4�,���6c�DU�Y�(�#�r��l��w�H��$�Y�}3��H,n�	�2O��t��j�I4����-��l�}��5٤�����W�l�ړR�ʞ)9��{��8�S*�¡� O�`@�zB"���2�����I�I�$�����\=���y�a�BQC�FB1Ev[}1ʨO)��b��-˭0�	� &�,����h��N�	{�K]MR��I唅b���9�� ��@�t�E�:���jmc��K������#9���4� O9���齵 +���~U��T�!���l�>�B҆[vk
��*�a!A�q��C���u^�qT�D �{=��6ec|<y�="���Z�՜�
[�F��1G"�b��=�3��7[I�FH}����e�ԣ��Uk�L�~�"nF㩛�X� �J!�{OM���x��� ��z�k ��^R��> �px�F�*8b�]�j���:�U6f5�a�J�6r��ă>�\�{J�l��5ĵ|u���Vgِ��Mk�_�.N)�
�����vǅ=��awvЙ4�S%ee-|��E�P�>p34��l�-���l(�G3�[��Ψ����`� ������H���X#I���ٌ���܂�TC$�&t�Gk��yR�}OY*=3l�D�|��Y��R�+z��(�w�f��IFjɑpY���a�J~�*Z�O4�Ł��[>h�L� �Z��~�I�'���! L+��[|	E 8}���t�a1�p��H���WQ��8s��"�،��0z:���5��
�}%x�`���L�ߍ��o���Z�Z@I��~z^ l��b�;��Y,�k�[���������P;⶘�)O�S��N���^��@�̋�6w��Z>Pp��|�ՙ�0�}�Q���Ԏ��V3>Q�5,p��[��%3�v��U_!�=d���,aLHi��*��6y��:��3�u�/�d�_�R�a&�+����H���,�>Vt���<@CB��B����g�+1��?u�?C���DU��P�T� H��@ٺlE)�@ӓ�
<I�H�ހ�F��:��?T�P�i�7@�b$�]��K�](v[	�钙~6	S�+��GQ.��w� ��x�m��@C��^�;J� ������
�QD)rt��މc��mZ�v�6/��g\���KS�&�Z�i���2�J:��˯xi��'υր�Qc2�=?�m@� �x.Ar$�:ܶ�D9�B���h�k�yAH2m�?�5h(�z�Ǩ�x��nܫ����.K7[��d�dF��?�R� �H��M�d�à��=3{�i@�y@� �u���&uš�5����&Ɠ�V�.�gL��lڻsV��h�(�N�*��R�û.�f�wG���SZS���.:�g�6�[�787F�}���' �"������RZo)��7p���ˈ?��B�ݗi����e�Xv�* r �1m�\H�����j�