��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���,���`�Q �����6�͍	),�6�md|_��n�x�"u������K �5owJh�E��qڑI9����%,%UEwf�x����;.�9��p3��,/�֤����"��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ�A�O�c9b��2���j�:��HA��?�\/��q�k��#W_�0����J杦�&���£mj��̟鬶�Pf�s5��q�Җh.�k�/��HJGS!]$�y�}�t+��`O�u�_|U�&x n��~���u^��'V��+�}Y}�� ���qϩ��*�Y�>sW���qF���Y��jJ�~�.-�KB̵�`X �!�����H�|)�@�o�5n �@Io�%L�}i��9��!���ز�����N��bG3���գΗ�Y�,G!�*IT���u�AC�/��1�؃z�Rj���r��־Jc�����Т�4�e.����KɃj 6*xL"m'~��`Ϥ0�R�A}�u��۟�_9^��-	cTM��D�w��[`��	��湟O'A�ē�_��cYl,�4�tw��E|�:�c, )F̋�"��6H����=��)�sDbwH����?�~�YKZ�UN�k|���}���-�$���TL������_��ƚ�����+(����`X��.k�E�O�BӉ��?��P�ɑ�x�׉�Mm�	���qt�[�}G tF�e\�#X��~]�SH0����?ip��_�f^��y�_Y��xFO�P�����8o�;V��I�6{BH���~1�{�:7*e�#�O��\�2C[FrM�Fh��ԗ�]M���6��k/��	͕�'��Q�k�@�`-h;O�x-�b1*K���W�(jjg�˭�  ��ϵ��zϗD�8<�n���G����
��g��U�Y�ӈ/Ov���7��Fq��p��jz�V|��Z���0�!��/��f�y>�Q�?�;�f�{ �e��+w��N�X�M���N��&J�Լ���b�E��ȇA�Yy��!@��óZ|�D����@C��,�����_��R�m�?�,����t%�&%�]�˚�v�l'��*�� �o/2+���X%�$l�X�@\���߆G���g�Fehan,(:�sQ2��L�al�54s6r'+��d;^<�E� _��8�������켟���ؾ��Q��k�e�+q���E
{�������G�"Z����1�Q�!I	ң�'`C�Y>�i1Sک�20e������o�^�,uw^!� 9��3� �ԭ��Cl���)�t��T_Y��Y�b߲Q�e��͒�t\X�_��3���5�j�V����Q���a�4�7��։5��6����J�=)�"VzI�}�������\�?�X��a��M���2�3���?5R�{M�N�'���b�<�Rz��?�!�vJ����:~(&匯�I$H�T�pT�=蹒�J��^kt��z͗�8ׁ��b��Rk9Ʋ׈e��+e�@�U��� �Q@�r��e%��'�M	q.w�(־���Z^��y�l������j��ݼĎAo=�)4,p�-�hQ�����tŎ0�-\���"�g��������P��҈9��>`+��q!�T��J#��\FH�I%�1���4B}J������W�t�$nw��Qo����&����}&H��ز���h}.4�x�9;�U�:��qK2 Ehdd�",B�~�x������l���7�/2P�B��D��^�� b��1	s�|�i��_�,ݨ���)��d5#�y���.��C�9�
wL(�H��f��A]K�����KwF ��Hl1=V[xD3�����I����MKY؆��>��P#ӡI�\�B|��*a$ /�����~��M�)rS(���M�������"%��X�x��WG�Q}��%���a��q�����(E��*��D-��{�����`\������Ԧ����s@؂�:���e0N�"�m�PR;�jmlD���/Igk��J���Ŵ�Ȁ�x0ܥ��<U5��W�ҜP����d�n\ob��j�S���n�
�����P�C��y-P�v�d�Ju΂��(  ��1�'|.z}HHL�����8���ؘI_K8Glf��IJ�$~
_|/~�<ק�mE�-�*�J6VY���z�W3��m.�xg�D���4���/���U��꺆��A�F�� ��laf%�~K��$����K�`L�-�"%���qq��Y~�{[�r�R�U��I��/�Y��FN�U�����%1C12�.����Q~\�rڳ�#�x��~�n�/x�`	�	�p[�b�ߕuzo�~�L�.�E��g��q�m5!�����?��
g�����bdzf�� tuB��ډ�����e���xw�?M,_�׃���ka��w��5N�@�c�J$��d�@{��w��-X*D�<��Ą�}��B����&P��Q;�xN�H�3��cɏT�> �ZLL����>��.�J0��)醳S�o��-h}|�sr��:3Q s�3Py[�Z�EW�?�_���Cz"������@L�w
7E�_��|�$�m�ZFe�׶rW�g�Z�H�^T���.,�vѸ.m匚��_	r��Ip0�.r�+(�S��F�YW+k�-!����~�)цj��Si�8���e�nO�����Ϊ>T�H���+N�=�jF�GM>�&`8�Bo .�f�;��%/� ��t(�`�Vh���Gy;������OG���;̸�%A'�a"tD��*Z Q��2�fq��F���<�3s����%k������)���g���&��Κ<���mәЍ�[�j���!	:X�da;��皓wW!4�=V�_������Df�t�,a��)�ź������u�UK��?1^���L"3�Ze6�����y���e��5�� J@T��7��x6�֊���Rr�+e��\���i%D�WW�g�)�y��H��k#?F��ޅ1WZ%5ˉ��hk���w~�vh�IS-�Cy.�ӊϾ�(�6ܯ�ɳ�K�6��hfe�aO"�3S�~��+�Ȗ�Ͳ�O��R� ��"�PI8J�΁%��39�Kݤ;ł��[7*�A!<�}o�p_�E�� �P!�{{�:����.��T�%��[��j�ds�0��Q��������\�0���&����w��6S}[�{v�Wa3��w�&+Ju�[9_�,��[k��V���+�b��%q�b=�cb(H��q��ѕ�;A��Z���8Ӡ�Гi|FO�<T�o�B�����{%ּ���?n�3L?�.���������C�N�<���Cv��IMT�1"�44e�I�l����=�z�g1e;����Lb�>�V.E��p���<-$H�>�G�e ���U��P��Zd�`����US����UhZ4����Y�;0����x�Ra�(<���;�<��T+Z�E�0A��䏼�:�aO��Y�)���X�K|D��Qv)��T;��ۋ��'^/�%�Y��5D�G���B�p$R�^Ա�}U�$������Vq;ϕ���c��m�X/�i��rL&]��Uc"�O?�+�g���7��d v;�5��n�@�)fN�RH�K��>�)�6�n�
��w U�e{c�ߟ���{eS��P�gya���X�)��tK�}�%zvDaƌL!k�m��E�#�(z��[44S��nc 3pa��_ �l��W%W�y�z���TΣiz�Z("�=���6����s��S����í�v��O#
9խ2��.�9A��zmׇ��[<�m9�����@���F>?�nO�
6�{��ߌ�9#[wIk��~� �;���]�T�O�g�^",+��z��ٷ��5~�V*A��'�e!9&fNs�)Y����Z��#�ă��]:����@�h�" ��3��v��z�5�ENǮ�hA�S#�h�
t>�[��������e��lD�'�1��{�F��-�=bVj����6G�$���L�>�0�IRxT��л&z@�)'�
b��<$q,�v,���]G<U��O�����8p��VX퀸����t�0�߃DY��ޓ�W�f�I#i��
z�~Z�*�JHe�Fqz��j�"�B��ՀV�-�e����U6Dɡ�~�.�����+�JAb��D"��qΜ|�	�"-�<|�]��y�b_�]�ko�Ig��ڛӺ�e�R�LvJ�q�u�jT�>�<L���U�W[�x�W��^�n �t�Ȋ"6V�
�B+��0MR>�5��¥��oܣ����P����X�<���u]վ��8ydB�3�q����
p�$8�4*I�`5���"!ZJTD\�����A@����@r�j����d�Չ�U�0��`IxK�g��@o��?a��-�Q'%�.rofR�n�ߦƜ��f@��L���7y}#�[���4�1W=�����:�P����h���a�"c���7Z�D��g2�<'���'�1uN��6�k�lW2>$J�?�Łb:^ʙ�r��2\�r���,��s���FX��7�7,|�a�)(��
�
.JG�ˇ�IU��b$e�F*�{���
�#겤�_�_1+9"�~mg��o�#4A���=V�/g6��.Mt���^����e���9t���f�L�/0��p�ĭG%�2������/x��o)]c� q�&cbDr�[�{Ae���J�&��Vj���:����\ �W��d�i��j�rv�nN�1Q�I�3
c�1�`�l!���W\��t!t�aH�V���8���m�`�s�x�
��X�2pn'�K�vQ1�2�p��������Qڤ<�ӵy��d��-b��7T�t4O��Y)��[	����.g<�$q�J!U������%ABS�ϟe.���0�љ�z�E1T��4�����{%���*��HO���r�W�a�y��*��}�f� =�~���$~z.�v��y��q�QmJ����m(��E:&���o��n{)��!I{W,N/>M��[Ţ��=#3������Ơw)>`pUl���[�;"�|n
�L	]{B�T�y��V��:؏��A@ω/{h�"��䒿+c���� ��9��`S�`L�Тv߄���s�v��ˈb���R��նܠ.�e�R� DWkf�#�D�{��05�2��ӆh���4ow7���؂������y� Ȯς6}�<��8�S8�Γ�o�00������'@��&B�%��ѧ�0��	�T�w��~��B~4�]T�[�?G����|�[��-���v7���LJ��ѣL��
UD��
K(��㠁��#����p�	�o�d')��_j{�5L₤#Yׄ���@1;N�X���I���
9����Y.�������zFS@&���{^������?�{D�Y&,�?��/���R�Q���s�G/x�u�{D�j���)Kl�~�YeFW��1��9 �莱���^������k�4�
�����K7��9��3ig[i~������Rb�9��Dc2A��<�I���	�a�<���:(��#���A|(+�
0\�f�XQAE������:l��R�?>ӴN_C��6N�BD� jc"�/��]�[���y_�z-�A��4]�L���l%FO�>��z�jl�鰚PO�R��M��j����>�����É���49U���ӳڕ8t�[j,����)T����03a����]�����E�T)a�WF���ӧ4J"b�)H�S�|M�ݍ�6�=����YfGY���m�c��偳�t�PT?_����O�?�FY�/ܥ_y�)[��1���$��c=&�jH��i���%ƠC�jtlx�&��ڍ�]��!��ܭG�?��v1dO|���� =�!�9�	�jO��B��"��Q�'0��R�~&�)��_^��cc���Om�nxׄ&5W���c�L�Ū\G�~X�q؎�F6[����˥9L���G��-�if/��y�5]�w�5�U5㏨eE<��?���y�&��3w%��r�/g�}�}�~d������]Ɔ���Go��Tk�%k�2�}ò�=�ɔ%����fN�z��S�:4�-���
�"�4/T���9�m`���1���������,ϫށ�)��m|��P`K��b�a�R�J�H�j�.�3�)'�0`�v��x{MG-���v�[+��on�%��Q�h�u'�ǿ^��X'	*�_|����z�
����MD���h,��h�4����0�Ŷ��Ww��P�C��!X��������&:*sjO�.̂P����AUױ�c*�@#���f���T�CWF6��i8$OI����
��ؔ(��G%�:�m�ҋ�Q����)�B	MQ%.JG��|��N�\/���9��t�ssm<m>6�Ҳ�
WZ���7_M|�]�5���/���RtC�����u�!^��儁B,At�9|��RzF��o	�
��N�]�r���n�m�s�� /"9f�g�W��-��"��Y���
-�tl{���g��qq�}۝� s�)E���3"@>����m�)�Y;p���C�l�.�F�elF|,�d���=s�['����&ZT�G|k0�,/�G`�۾�W|Ro����Uթ�����X�%E��~�4��;�1:�"�r�Px@���<sOxZ��@��cf�&�m�0Ҙ��Gμ(��w�x��c9�E��L��u�j��m��/�ө�$�9�G|џ����	m�3��&M�#�y\�g�A�$�<�2Y��x>CRFt��5�����0����tm���I�%����0�-��������8� �c�*��Dd}>s���ڥ,3ɃzP���U����%Oy6CÛ�
Iްi��Ӕ���'���R'<Y�ߒ�����$�� $�H�ܴ�:�I�6ڳB�ȋ���'�.=;9<�Z['�x/[��Z�aˠ���$a��[�HȞ���-�V���W����4-̊L���n�*����ށ
;sv�TYuU�;Y%�:lc���5��1͈�n�.tR�C(6f��uAغ��Q?�]#,��U��l��^�m��h��j���=><�Q�[�ri�N�=�M�����*'�O�(��:Z�nW�f������G���q�e�k�P�
�MD���!f]L��ڸ	q}���i%o�0\N�c�uG�ٔ}:_�4	
�n�x
��]��I�jc�J�t���x�a����{��%f�����í�r�W�������_�Z�ӖF��J���(��7�0���)x<�f��q�\�Z%�1I�BY� ]������{߽8<FZBلj�	9��*.uo��)z����e,{m�Zc<|�����u�c�> 3^���q�K� 4s���T��L[�ra����H��g�k������v�q@Z��.�Av�U�I2����/�f�9#C7y���;p�o,.�k��%�?���5�M�g���'|���tߞ~<�$�D�>v�������	��.���U����8^�b����Vv���~���@�t����9��������m���g0���#���1�퓰�O ����f��:��u��/z�D�F�C0n|��)�������z�H��P�ߦ

����B�&��d�L<�˵������,C�]���g�vk����2�0h4}�p�zTā���:
�����	��g����qx0���|Y]�:+K�K�*^M�����.��m;��s��~]7�.�oi��!��~��|ꁎ[k���O2�j����溼�/����H���~Ҽ��<1 3�qDv��LZ�b~�M���ku�B����5�;< �w��~J9 T���j:���`Y%�]c%:rJܜ��U6%FI85�s#���S��<�I��4�e{���Aᒻ�ZW2V�vÁ�e$�n�B�\l%=��q��2��S�K��\>�jm��;q�&�ZS=�c�z���(��Bi�P�E�B&(d��v'�aPK����>p�����j��}���i�)g�13�W�I�U�D�b�T�~~�PE/`���C`����ZgZ1�_�j�-��3x�������r�:Z}��L̙o������H����-	�"	�۲dx�M��CvZ�������X��:a�b`����|��l���]y�����p]S���9�k_�_¬H��Mχ���9
�:A���p�4��,O=�?
����7����4�i=��c�U0�OC^|�!h�l�Ғ�v����ǩY2�����e�)݅��֐��=��2�kF; ��)��g`�z.���S���W,��E��J����[q�;Xd��B����'g�9#ou��u��q�qw
(�0�(��ـu��:��$]o^B�-�|J�i5?�@�~H�n�\�'�>Ԓ3�C=�?�\�#��� U]�I��o���7�]yG�/����H�i)��Х�B��(�_�Y��XH�5v��x���H? ��s�?гY/�S�Ɍ[�<®��1͚̾��d����R�̋Z�2����o�r�aHfI��|<����,�ڲo�@��4�/3����rӿ��6���6]+�����@�~��	��nɱW9��	�C�U�6(��7==B�dp�`�I�'��i�O���Q�|��81���rO�W7ƕ=5��P#�4���(�{ᰓAB'�H�Q��{Bצnr��)xy�Ҷ��4P�q�����I���L$u�����L��7�'���?j�ƽ�/[��>�F~�/H�q�4��(_��Cc�>��rV�Pܱ�O�����"�����8�t1�h����Ro�fJ�}�h=�jҁ�E[x��������KJ�?� ���%�@��b󜇎[Է�UVk��O���r[�0�Ga.jٸ�����.�����0��zS�:d3��u�?��g7�<D�_kh
u �Һh���O�t��>���v�i���8P���y�lM��o'7I����\��= F��Sxo�Qb KD[�΅���oJ�#����9K`�+Xށ��蚩y�Ҥّ[:leyra,�����k��eQ/մ?��#|�c����"��-�8��ctC���i�-��o<`�XP�v�/gC^F�O�Ԏ�v�'O#�D�rm�/6����;8�DU���,-���k�d�:���͕�T*I8�/��o�W)������$Ot>�A{���<��� �<��'l*U��g�f+o(氹wE���lPp�>�΂�]g	��5��7��Ճ?C����C�K���C�i9o��%H�����Np����a����iY?���������e|y�'�����E��vy�EnR�� G�3wM������u�,麰F��h<�W�QJ�pr$��"��އD5���x,O1�*�3q��
��[��*N)�x��zM�$əpPv�(j�v�M�R,)l{����._B��!k!�v�a(�\�t)�ѲO���v��u�H�}k���[��N�k	������զ�D�l&��;8��h�uݓ /7OwF-�q-7%2�0R���0	kd����\dx��_��@Ȃ���&���頜�)�G�Q�\t	.k^�1��]?�M�]Qou���+Ѹb4�f���TYJ��][g	� ��ˌ­�a�
��#�p"�u3�-�;�p�j��d��eV�c�~z�e�;o�}l�2L�<4^3��ٹ�:��Hߡc��U��я�%��m����غ)�T�2��������t��6X��8��'e�[�8}�bw�l�,��B�	i�)زP�=:�B�-ˉ��:PZ%�T`��Ʋ;xG�������0I�a��u�ʗ0��7|j`�/%Deph��$s	o��ûю^#v�`s\�WL��:��� ��l$���o&o��yx�cgl�(�L�����8K�1qM=�>4�!���en )䰞G����c��b�Kc��輙�ΰn}�"����6OE��%�Ў�r�`&H�8i[�IWK�T�yu&+|�?{��� �i�{�և1�dF��b��8�wX�Ԏ6TfFQ0��P�=I��h2b��$��Q��O�GQ�#���T�/+'W�
n�OP�E?�M������!�|�4��>��R��H�ˏ�(뙚��㠤�G�N���R��%|�+b�V�KL߭r��Ɗ���s�%�P+
�4m@=,ա5(m=�2��+]d,&�� �Bc��4���d��l�bI��,�]�f`@���-�-KS�t����p��{s�sa��2���ij:N/jn?��5+�Z���U?ر:7́��qoJ[��l�b����W���"r�3�X��}Pߔ�]��)�}�O�;��LMnHl�{�*�vafS<�+��p�z[G
�{�}f��E=��,=}�ow��'/����Bm=�X��'�쾔�]��5���ŘF��(J*ChF\���^��� 0m��y-v$l3x!Иrԃ X��Z�Y�J�>�:P�H��+�l�A��}L���l�#ljz)�~!؝��7�QL�菬
༄t�7����֓�6g���f��aI&vJ7�T�8�bc�1}�v?�8���_��)@Z��lx\���R~Z�y㪋�A�)4ƢF\���w�𚗽�Iy�.�j��d�`��̘+*��A��4��RJH�sM���*:���9�(/e ��[�Ik�zQ��"��}�}q�� e��u�}��K��(0�F��'s�)��2<�����=�����a�	!�����\w���}��-,��i�C�Q"6��}�&lS��)��ߥ֚��F(p�Ap�	q�x8�J���G�Ǘ��X���@���Zo�Ӓ��jJ��Ϊ�)e��w�"L�����ϰ[���d�/橘x�
���)��K{��dnFX�pQ�2��0~�%�!4�]i���9�I(��^���3[��9t��4�D?�&C9��`��D�+a��L�U)�!�����H�����f�2d:��.C�Bf!�D5����N
>�$�GJ0[�rçO@i���RY۫��9,\��;V SD�J�KY��=ck��C��������QS�j��3:��f�ո��^����o���<w�Β�+��s���ãc~����t��8h�����$`� �s%���HK����"��W�ɺ��� ������a�^�Y�ڏ��}g��Ϧ�n�|���⏑�It`�@~�EU�0�̪u�d��^gV��2�F�`rE$@Bԟ@�?�