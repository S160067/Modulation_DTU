��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����>�S��fI#�l7x%���$or�#�6�y���N�i� �D��f(�:eǊ�` ��S���^�mBƱYjA���v�0��kh������#�v�(#W��ux��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>c��mW���rJ(���/	���~J`2F�x���4W�0V�y��l]��X���8D�G$�ۻ��c��rk�E8o��W��z�����O�Q�F��?-_�䰹��Ny����o��:���l�,�:^�G���G��ta�`����k�s�|��8��Z���\�0��c"�:t#|% 3�J�o ��H�NS@>{z@�4�>ÿ_1B_�V���!�_�mXI��rM׃�4>$Z����cg�5x��H7��P�-̗&�����!)����sFj
rjE��E�q�[l�]_k�(,��v�:��^�g|?�O�`�亨��(h�^�;OS+ȥ��7>v�g���w�k�U@�x�tSa�ŝHXD�`��a�X:�� ��u�Xb�^��*�g�x�"����/޾��"�a[�Y�rsϠ�`\����vܨ
��G�<Bd�c	»���뙻��'uH|rh�~����\������Q2 [��<�~�/��/?*�D�shW���Yf�-ğ2��Ff�v)_y4��߱��XϜ�5գa��j�9��xn�uz�V�%�2ruZ_C��ҜO�Y/��a3Su������-�KH(ɤl�\Y��1 d=��QX���1*�	�|q24�]�藘�/t�k���7�,z�'ݨ!���� Ȣ�������ΎnP�&+�dZ���z��A�:�V�����w���le=)#Ҕ�95$��]�XK��3�p'�Q$�@�ًq)GgJ^�
���J��WH�wTvo]�I���0�@�}�¥�S��L���t���[��}:���b�g�ɽ��%H����ZMt�>���:�'�R�[jPD�� �ۆ�0����[v2'bQ���)�5�An���s��δ������D%�WyR|e)�ح�+��@G�^ zf�\�h�k�	zm��ǿ0J6�h;�1���-{���3���>�yT՘"�@��>�M)��S�y�P
NBT�x ���	�C��^�*�W���
�K[a����9��}aj�5�9�(�#t�U��#RgVU�I?�y>s±g��)�\m���+ok����XJ�hw����g��;FsH���zO�{�z��������"	��$� ׈���PX�����}[R�f�~�@�"������b%�c�!M����u���c�#A����27��=�{��o*��:�?����'�oJtԆm'�+��w���颊�M��L��j\��7R��^�p5�{�'V�Ĉ�\�N�� �z?�5��e1���%����V'��MD�3?/'V�e�����k���֏>�Ir=�����,��X���M�r��`�
\@�fn��A���h���*�3m�v���>�i�b���#������X��*c��4u���4�օ)I�*{��X�����as~�;�~ ��I7�L�
�Ȣ,X���b+I�*VH�� T��.#y�T�:��5��(��Ng4)�4�.�U�l�Ϗ�͉W��?	9�9	]��Ȫlo������:~���pMl0\�����S���G�`�8E��\�^R�P��zS3�%�q�jU*yq�aw/�a�+g�!m.������*�cu����Qp�-꣊g�%���_����	⫐�e�Д�-:oYGh�ձJ���A�cU����Zt`U��@+�6\9��/|�
� ���?&B�^�bL/�@�����Zt�]���kf֗Ջ�*q�,w.HC�Gv5����p�^���쓳RL���ܤC���R��O�dX�{ 4,��S���O�|/�\4�j�aݟ�D���(����/���f��5JU�Ub��ݷ�T�N�6�'I��R�e�@�!DW��VeR6�ŏ"(�"��s|o��S����}�a���}��&f���[�|������|��6��d90���>�>a�ّfAօC�x�V`[z�+���5�u��`p��B-����<&ư9٤|�m$wj-!#�?H'���E��-|Wdo��N���ϵnr��\�g�~�٥{M��d�3Q��~AV,�t�:\�]�����(�#z*�������鴑���l^_󀬪]A	�zF3� V���[�Ȗ�(��s�w�i�(�[�֗u*�kR�k^���t����Y�G����906��
���r>�����9���J^a,�6�ZІH��T卶�,J�R[RGc$��0���_�I���B���n����le5�3���1�/3�}���@�M3� /�z����64O�a��O��ܹ��~a&�os&����b�mBEC�a�����8U"H,jr���bw���9�k{���'�
��qZ�^K�}o_{ C�A�������pt�%�CbF��'�:��VȂN�]���݊T�0oB�'��5H���q������Q��y?~%�^����ԍ^֫�Q
;�<���5���k S�:0}�t	�=󖇎�����'�'���]�45
��@��|ѣT0DF��vZa.p��_�j�h��>3L�"nɃЖ"ɦ'�	���d�P��2�6!0����`rSLM���I�*�_QO��tTag%]�L+���ǝ5�ߌ{��&�[K	�L����[ukF�aR�6���h�c�W�� �	��V�8<�߳��P����Y���:!�	s����2���)���l���:��s�5�L2Ĵ�i�/x�������*O��n��]�q<!��!w��f�&N܅�V����{ܜ꟟�w;�nni����U���<u�� "�?�NTip
����sj�?�>o����reCY����[A������T��r�>�X�Tzp@��E�Q>5��Mb��wM���Lk���^vh�HK��l�8o��Xf��7�EN/��Ӱ��+kj���R\�Z�.�_p�!�(Sz!����>?:�0~�2�6/|ђ���u� �(M��pns �u%s� �-ʤ�l[�����Ϣ+1d�����2������U�q<?T<K����#K��Se�b��Ϯ�q�6�xw���M��lmp7�F9E�t���-��U�bЕ�������tK'�Hը��GޒUe2-�F�]����Y.y�v�^�\�_����;�Ὦ�(ª�W	�D��t4@���u����֏�`Z!����ڻ��Z�G>�TUu؎@���ў^�k-e`C��9H����ފ(����s���n��ys�D!��vб���.&*5��e�P��C��x�A�(/�\�j������w-�h��n&��F���Q�"['��-���dB����ʥ=>�m���}�sV����RDH%	��%��7t�Ɓw�iKi2�p��?ZH�c�u�3��oKC�