��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����>�S��fI#�l7x%���$or�#�6�y���N�i� �D��f(�:eǊ�` ��S���^�mBƱYjA���v�0��kh������#�v�(#W��ux��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^���y��Z��(&�ς��%2�����1X���N��x}_�Rd�`/�-����"�'�S't�+"mRUp�J����9M��}n�a���`����*F�	���w�4�bu�lw�6.0p9Cb��q�\�T?�/���෰�=�0�lcy{{/M�	:[D���ua��yyѼL�B\�n%�o��Fj���_eOfXY��7dB�r0��o1�2� �1#�g�,�w��|6�x���~���) }���*�0}E�C������z�/�P�#t��[�In�+A���g1�뚍u��dԹAT���W:4��ټ�e�Yӥq�h�+��<V��<aQ\������:\ㅎ���.~�<*����.���Fs��2�i���6z���KQ%��B��&c�!�D����:M�O!�"х�G�ظ,x���	�F̈́�tV�vS���]�������65Z����˟Y ��&(���rLo����X��FK�M���n���+�(�����#������{ρy
���Q���+Qr1V`����{�\~�^�d�c�b���9r�°"���b��*i����% ����0l�h��.l+�S��AjkF��O�m'c��.6@z�"�L���G����d�`u�e	n[�`J����.�z��"k�6cG��+^;~�n܄�r?�gT�F�Z�H����i�����1Ð9uY���{���Z��?���t����ѥ��p�&��u)��C��J�]�z��ۈQ���|V�@K�b��h�HR���hW�K�:��A����%��kC��=�~����\B���Z�{�j��vJ��W�1�e�I�I�����4���c�����O{�T���e�@�e�^��Ї
�/R�w�`���JV��i��	�]�ۥ�W'�@���!k�Y�o�s�v!���f���Z���`G�5��H��vD0kDkʛ�D=F��\�B��d�q��6��������U�{�����:�Β�8��؀Q��ttr�P;�辰eW8�����������bS�Ѣ��*�����"����6��
�y,���n���9��n�}��O���醰gT��v�!b�n��v�k�S�B����Yt�]X\��A��P��� ɷ�H�/TU~��
Qi*m&�g1N��:�&RR��=�U��������d�ܣ��z���y���t��J��y�[}#A|L��"6�R��R�1��uC_
�V3i^u�=Q��Hs��t�$�B"Y��Bݩ5�����Xb
���Ơ��K�zB�l[$Nvi�!G�	�h!h��B�皙�L�ν��^�؎"�����M$["�סD�	�E�LF�j�7�jx�}Ŀ�m�KE�%�J
�	ů�yVL2	dn�-$�����9d�5խ�|)��2���aN���_Ni����k��E9I�&"t�I ��~��f��=qk�;�_tƀ�sr�	���B����u�|�E��h�}a[�y�;����|�ͱ��W|�9�fj.8�d�������ko�
�Z$]�%���Z�O }��ަ �˅|�%��L��"�O�ѯlE�"
c-���.��kB?)�_�\�����ؐ@��{[��v� d�( �"�/t��v�-�t,7��<DAŇ+b1l	���q.��#��V� ��w�U?����X��X0�',}O+c��*��5�[@���N j�h(�a&�5[
)�8%f�D�J�P%�O�����U�GA�&O��'2����$�D�ciO���ļk�~o;[��t�&Vؒ8���vxȨu�|��mf�R���Cx|�@t��̹��O�n	.-e�[d�L���Q����������?ɜ�/Me�T��*��3+�9:�"�t�/��a�-�\VZw�#�0��;��(�|��$�y�³Ue| J��'nhJ�#"�fȸ�&�(�_�1����IP��_F��7�\���8x�ׅK��̽�Q��]FP����j6~"��@����Au�|r~��ϱD�)���E��|a��={��:g�-�z��̷���i��w�S%+�����JPZ��Z(�7KvwO�����H^�jK	}�1�hf"��g,���`	1e�� E���s�ȭ]�ݚC�B99`��C�f�s�^"V6�o'L�X7Yau]������"V�*<��GF34��Q�9��g_�#˻ot��d0��i���an!�H������]w��9l�T�m[��/z]���E���+썄�Q�4��B��H�aĨ��k���oz�4���&4� ��OzV�c����K����M��S!���}�l�`�d��(���ĤK�N�qٓm&�2�(�1|$�/�I�i>B�ޓFvonP�Kj~tZn�D�s�o��x�| �t�E;@�!Q�`[����Q��IY��`s]!P2�	f�f��㠷��7a�%`��?F6�'�x>p7Ǝl}X���Z�z-T4i���2W�ӄg��q����_������S�pn�0#	)��V��Lp�(k�'�Q���X���z�n%x�E��ݻ�Z�������=W��y=�]J����nW�����Z�C#F��q�n����$q�T�xF�5sd�������D][�D犧�yg�[���$�������9ޮ�� ѻS
]����d����Lπ\�X�	y�̢XӠerW����*GE�kS����^������%-�C�κ֟4��4�3`�y.���X��T���NDIq���ޛ�vF���m79�;x����c=���hN����frQ_gM��R
Cc4����)��򗭤U9oa�О�u��`���Z6]-��z�Z��s�{b7�=��8w��KÇ ��8�Q'А4�p!���Hϲb���u ��mh`��n�FC@�ϟ����yޜ�e�h��c���,_h�5�����p�`��&�*
>-�C�.��R}ǫ�e�À��	�#�#ͤ�<;��r�ժf0��a�c7+�3"����qX~���}�{��kG(tSӖK���1Y?O9d��`Ͻ#�~s��v\+o$��f[���R�L�ۄ�M�h"��� ���4�i�U#)t�>[����3�hCu���&0to.N��߄��ѷ��������f��yS�8�О�D��� c-�H}�7��2��#�,�T��Ǯ~�J�����k�y}�@�+�(=�k�Tl��Y2BeCZarj�G�Q�X}�С�����1�e��~��y�[=�3�g!�:`�Cw��hgq�~��Iyb0+�ְ��<�K�t�(R"_�Ż����/���j}�ɗ&~�	,4g��p^�~����>���|;/������� $
z�Л�!:��;:,�M� �s �����EY�C������kV!9��z��zO\{r��bg�ɷ��
���yw4��m�2p��W�٤P/�[��j��p�>;���]Mz��x�2=������ 9�����-�KL�z�O���L�9f:�T�k��%\�>?�w��iYk� ����^K��T��Pw��p �=F�����j]?���0^<�*���X}�o���iNmx�Iͯ����f�ܿ���ҋ�T"d*��/t��G�s�)iLI���Ƌ\���#�G;���ɾ�+q�.���������+������D��p&��@�	����� M"<�p�6z�tܔ<�צ̡�^/���'C�NU���Y�B)����`�p� �*�k��BY����{;%���{�{�1Z�o_e����ݎ9j�5�;�)�~�ߌ
1� l&�33O~�"N�����OFxU��U
(U��n�:���dZ�R�����	y}J�(,��@:�?@�����੸�Gx=^yç�dE��H��f���~�l�Bp���
_8�{��f�_�}N���B_E��D�� �u��1?ʖFPXot�� ψM��ˬ�L��0���P#Y�;f>�M˼4W�O��'٫����!�fP�WP���W�o�S�wq���f�p���x�ԝYF�����m��a�:��i8t��@N,�4�>d�`�W�8����ϯ�a�0t���+`{3*�����$�뗇D�GV�QR��@��"X�uZ��"�	|���`�!��:���q#2eVJ��U�,>�v�T������v��I||�:����Xa�g.`2#^,HaR9�ZA�X#�Kͨ��ƞ����<��T�}]ȓ!��,��	[��I�%��>���ff	�W:�4�?"�����DWc��5'h��|�1�~.e��ڕ]>g�TC��[R�Ҋ�;0]��؃Z]��#�D3]ٵ,c3�C2c�\ȃćr6�;JDy,kb��:!<^���\Ú��RwaV��Nw	��>�x�I� 0�Hyɪ3�g)kr	�'$��,A�%l�僽�Q\�Aʍ���<$�%bX�溻"���u����B�׾�S%E&�dU5�
Қ�T�J�g�	\'l"�����qv��'R��-���I�0�d��򙦣U]32ݬh�@@�[�h�W�
�Ֆ���f,Z-��^g������������ﺊ������lPiy8��y{�)�YK�Q��D+ߑK�ڍ��ؠQBGVb�m�RB�mi�?Sɓ�r��dRυs('h�̶���Q�0�I�����H���7��C~�2p\qJ�����ƔA�ͭ���.W=�k�{�w%��:-3�znO�Nq�bQৱb���(�퉽2v���tS��uNT{!�����n��E��4���� c��B�0,ya�	��<��hܵ�Q��KR����S��&�K�j��ZjL�_DQ�޲TO��
���iĪ�K�7��~�C"4�k
xXs>�U����`���:�. ' u�~�V���~��Am+���\鯞�6k;Vބ�oc��h�w�Դ��y��r,�1���6J�بF�w.���Q+h4m�v?ŋ`[�]6>�^9��I��Yo�f��{y���|S�?xdw�0�$��\�ASW��mS�c�q�V*�ϹP^��<��4���DCۢe�-|��񦮞K�P�d�(z���G%v�.���I�M��<9ˬ~ɝR���}EV������8M�VfO1<��5Dת��~&���X<�r]��<?$g�{�T�?��׵��s�rx|���?��f���9�� �67?F�t�rT/��x���Nj�0Ă���LzS\�ڣ�Yf�m�.�d��S�i�KZ����  ���;M�}�='��u��=�l�k�GQp!��A�`|t3�E|���#f�R�gTl+SPf �_��&/u��G�|�^���m���}��&}���j��c����ԩ�M�W���iC�����U0h��R&"4����zH3{8����1�b
���=��Oֵ$�b�g��M(uC鼪v����ϸ�z�p�@[�«���`��R��>�lP>���a5����ڔu|��Z������Bsmkk堆݂�R���'�r,��V#��-IR7S)C���H���]Q��R���x�r��s�uV�u뺐�����cHl@)��h�����(���i7$�Wߐ�\zZx\q����V�S%I`�h�߃[W[b6�ͽ�e�`�f_#6{��/���H�0���ѽ��7���!)��h��$�p�Rg�J(յf�����7d���"����ۃ#ρ�b+7iY�g����T&�Ƕ�,$���s�I`�Va�Ȝzр���� ��\K��l��D8���c{���D"�&�hV��!��D��Ԯ���T�ITZ�	�@('-�;�d�"���]"�a��Y�ɤ��MQ��P�f��h�unk��h>1������U���d�bl�aV����c�6}`gt�˼`��K�+x�2��cЯ�R��G-��z�	�\ԁ�+����c�;�h)	OY��r_d��N�d�+�1vs8��'7?�En`�?bl¦)|y__�n�p,�j9��R߇x0 �F��X��q*��
94����*ᡉ�:q=v��p{ �;�81,�Z���t����eز�P^���|3��"�x�hM�/�7mW|ʮ�Wc�?�8(ۃ�stfr��D#�"Jt���x�jv-�Y�4S���x����ϳ���&�[��w��,R��Ν�C��w�8����A�ӝ���3�V�0"Fu�
M����%�l���SB֭7ƀY֡���E�mkb��0^���R�GPd�!'�Q�?u*Q��Nk�=G��4,�6a$� I����R��9��Lp�E�4��y�I���DUSS� �aw�~t�	J�38���η��.�q��,ǂvI4:9/�W�'m/yF}S;)��eF6�`a�[:��ٍ}�v!9x\�}�Ab����օ��{��[�<��o,�Y+W �fȝ��)]Y9�t�Ԥ�X٢
�e�Rw��Kb �S����o�%��Z�
�%�lŦ����f1�,������!�[4L�my�X����MER�ί�i��޹�0���[%���!%�?˂�D��䐅d���Ǎ����?-����?F�7�i4AqyU'�nT�1I����,���Сs?�.��ԎP�r�r�n�(&��������fk}H��}��5"��A���D���M���ӂ��"��͋'���V[+��ük50�i����a�_� g�����\�Z��0�=���3{\�h�\��ľ�n#{�ؑ�zfB	Jʥ)}_H�Te����z�y���2�[ð��糖u�̪Fv#Q�`�J=�d��]�����XE:�8ƭ��ʎ7
�l\��&�=�����A���Է���S�`�%Q���2�W��_hVY�4�K1̪����Vo��e&y�0kUw ���ͪ��15-f�,.H�;h�*�7���؈e��L�ym���fG�Q�WLSdZ�3`	[�Rԟ�Ձ��& �&}���P����{�EEO9�WrM-E�\�q_�TӱX���(�?�ʗ�v//��L���	�㼞d�'%�2���<�g�*���w&g����Tu�Z�Nͺ.�8?MbW�<�����E��x�Nc��T-����r��M��pa?�2�X�'�ZξP�"$,��H��B�jˡ
Q/m���"�cH�hB1ݍ��Ȼ�O���H�x�7�T�8��>��1�).�q�`!� ��<�����N���S�B"�w^�d��l����~$YE��DtJ\�=�[K/N�CK-��Sy=z��~�B�b�Q�a��,o�^@��_G�Um���3�����1�g��߰h8��=����CA��o��8�_
W�:�
���Bc2t��c�������Ĳ����@��cH���g���@�n�u�p� �P�Y �YD��.��֤T`(�7%�IM�����}��̿�>���`�A��Ppˀ0t�
�X|3�M� �R-��Q:��6�m�Hw:h�L���3A<���*�O����n�iۺ��rg�s-p�䚎��{2|E�>�]�e��Nؐ\::��wM�p!;߿v���8�H�������<��h4k�+���N5����O�?�RXO�"��;�3u��SE9ʥ��@��Sk`�;��;O��~��[��]� �����e͗CESt���#S��b�����Al���r�9,=�^�17�h'��
�p8�X��̝Puh����p�5Ѥ*O^�@��=�];��z���v�"�Q����O;�7t��%z%��%�=y]�LAK��aGbC��V��h�������r��ˢ�e�ݩ�'�@�����y��ah�h*���}��t|�l	�v�A����^f���>ݯ�U>I�����]�y��XE�^��e�xiF���Aa��k���Y�|y�K��*����߳Sl�#�r��|9�qU6���e���mL�>�T?��9�F8�`�[k�ݽF���{�r�oZ`�3�<d>�
���UT���Y���|�sd��b0��Q�!�L���������n�g��y�fd!�x�摄�̃�/�k�� �Q�l4�ܣh���T0<
�(&��E'��^����D�;�ӿ�t�m�+�H�HEFE	�i+�q�_t��S*���i��;TWN�?:��"�r𫚀�ɲT�6���B�O��\Y��I���u��[ʶi������X�a�}�D��~[#w������'M����R��ɏ��7j����0/�r�Lح�v�����\�X=O'����Ug^�.�H]?v�D�k~�|nlsݫ�_4�@�o6�W�\��e��8����c�;�����	�oc��u
sVդU;?j�}�$
2)wYˣ�
KYk�Cu�RY�-¯���\N��L�����Be��w��������ｫ�Rch�Gҏ�':��ŀZ���+�)D���+P|�D�����37,�%WD�%{�f�jb�]-��C�A޴E2����ʭ���� \UJd�o�#��O���5��T����+e��w.I!�N�/�H1��������EǆIc2�����|�9K��^D���@��֏�{��ؙ�/͇��YSK*�{�Z��bxh�>u�=���o7}ԺM��ӫJ����k�`�0��g\��O�G�g=�5=d0�:p�x՗��n��b�^k�N"������9�µ8��H��~5��ݕ�y,G�Q(�.�c�Xjk�|�7P6dS���5OY��v�=H���c˴	ܦ���ip�.��u�Ʀ��|�	~��{[����H��3�\}���(^Mk���A����
�$�W�t�\o�=Cc��Xg�s�:�+�k�K�]F��r^��mH`F����e:�
-�t��{f�P�� ����qp�c�7ҕ�A��BG�=$,��m����tq��5֮��+$��W@Ԇ�9�*�#��&�INo���~��l�CB�~O<?��S>ϐ��ry�bH�VJ���������G�{[�E'N8ݾ����Њ�8�l
Bw��+��zI�:��l����|f��p�3��L�]�?�ݙ��l�@=��?��TdQ�<��LWr�s���s�އ>9ҳ$C��E��"RKZ��EK�)�k�b�8�I�N�`�i�驖��2@�GV����P��L~�N?��P���2#D��شH;�WuܭN��,��gK����I�7��i��Ŕ9N��?�^�.ρ<d���8����g4!A�#3ʀ7�lP�ι<��T��u�����{�d�����sk��-ڐ�|�����)�7�C={C0�U�	�1S��<�w.��Q��s��ω��%;�mW$ۘ��ێF�!(-bj~�YF�����T�c\�i�5���Z:�Z��$��[���?M-�&�@�_�V����g�h`#P�,�\I�g&��KG�;G���BVh|?�ѽ0����@	әH =T�����W���Z����<��j�OS�� a�I��<4xs�y�/y[�n�{�@I�ћ�D�����.a����uc�����\�r��oʱ�y�X�$g�&@餛�QD�tb[Ǧ�����M;uD��^�Ӹ8$�ey�n�TR��dx�d
��vu�嬖"H��gw�;Kc��
����s�K��j���>�.�oz1	?�D�k�5�T�D��mu��
w�p��+��M�"�=;d��,���̓��#�Nbm�C�M���?:Gr��qM�,3���A����f�EZ�8��)��:g��8��9j{�n|�M0�C�d�y7A
B&×��SFV���j)�_��ED���/�[&-h�2�����3��������C(����5�!	#K���<@ p�aȾ�@���)bv���Ì��r��JA�������S�syGzR1�E��|�1��F���,hGr�b��U����rV� Q���L��4�}<\�{vqg���䋲U٪�jOD��Y��!U�Gx2׳�K��ל8z��2�.&���Z�Y��f�k��k�b@�������(��`��C ��n�Nj���&4g����70l�O���7�)!!pc�|oٰt����$�[_���_��c�(�L(/E{�Hl�xB~;El]!2`	7��$���1�	�e%XeY�N�(g�T#��:~ �އ�:KU���f	 
5�q #\�ߦ>�Ŕ�j,��?Kex�8�P���\���~
�X�'�wF��Տc���,"�N��V��#Fay�!^5ǣ�v��Tj^�<���Ƣ.�F�\����>���|�e���h�j��2c���@���@��BW7���$���d���M����S��5��i!����t K�{����|��Wc���ɜuC�q���:0�������p+��SF�ܬ���9�@j��D�V��YpX/���:Y��UM6kp�αy<�pc:Bk�k��BX&�5c�;9w�Y������߼�H�}t2e���L��K�W
i'e}F��+�4{]����W���T���Fo��T
����a�C�m���*}��'%x���$A��*��;S��!�v����ڴ����>��,�ۇ:e�ZmQ�h�����7�t/m.w�#�@$�c��ĝK_�/��O�E+��$��� [�%{��_��*���\wy�ļR�{UaM�Â[��`T�\�̺��Ei�]��{|�ʷ�:�6����L*���`��~LS�Kg�mo��EX��c��ȵu5Z¥d�h��F���M�Z������3���_!(bA��L�=�}�&K������ⵙ�Z�%�	}�V���(c9����>L�:�8�c���C���e�)�D�M�_PYu���)��pEe�y<�Z�W�aɪ���P0 �-5*+������Z���2;LqсG�aջ�j!]'����`�Z���������k���M�C�J�mo��@[
q�g�%@��ڮ��cb5jy�z
��rJyQ�.���� |���=�մ�| 
��i�=��sK)r���TE��q%z�o;�Hy��NM/hԴ���ә�jA��_O�D8E� �����y���������")��Fa�:y��u~�e��ᢦ���c�9�n�>����Q�ᗹh�R_����U�Z"�\s_/^���ymB��;K�7������6�x�;�t/��@?��N/�f܆����=��d %�������`����(���0��(��2�K!��1���QS$1��a����;>ޕ ���Zc>
D'9Oĥ"|��.s�����lSP
��'%mdYڵ8gӹKL�_��NB�ˌ�2�ǧJ�̅��:&�MRnRa�j�H��9Ϻ��6�t�d>_�})���O��c*=vo�;
(s�Q*ƹ�M%,�YM�� �o��T�t��]������v#�� n@R�M���-��ZA��a���XW���R5Q��y��q��	�5'~'+�^Bs���1�V>��'	#���l`N�X���x�Y�Q�����)o!hH6V���G:�d����N�)(�g<+���o����i9Sfz��>@s�:8��=6����0��PA�f��.����uH_�7��I'$����6��O�R�[�߭,E690׌�:����e��O:6�n_L�D"�K���*Z'��IK�p�Ąç�d���w�/f���i���ėop9��HC�W�^�`�ה�1T��TI���٣e��m���bTI�8�>F6�p�@[�27{o���P����
S�'�^c�Ԩ'�!�邂��p�ǁ�E���S"va�1�}����c^�mg�l4O�z,_�����@���5�@h� a�ܔ�J�\ix���t�i�����JJSƮ a�!���G��y���0!?���0�{���ʹ�C��BA�z�/���h��ī,}dřg���5\�������X�+:b���'�3J��]�_�q3�y�ۥ��S�� �_���FR{�	�OlL�C��zcT���A3����=.��y���AZkC@���.�
�O�-����b�#.����)��) V�ϐ����ƺ��`SA��d#:������l�>w��MCS�x��n��X ���>�E�*#Y�G0����}_�;hH�s^Bt]�ҐQ�@'��_�_N����7�>
�<͹��zwy9i9EYt���[���/����r1��" q7���~!���>���[�����O�����I:�!G���ϲ�l$�6�44�ҨW�Lܶ�O��`Wi8���#���]�mu�E~�iD2ϸ���߿ko�y������84�ޅ�=X����+b�PE��`��8҃�Wͪ��6N��{��ʜ�3��^v%k�*��Mc0lCU�r�F�vvg7c�`-11��;�����A�u*<x�v�W��B���48W���+���OV�d�"�i�	�xG���4
ȵ;�2���� �Rܗ{C*rO9C����o�Y܋Z+�T��_�M7t�=�v��5�gp��������\ޑ�G���qj,��������`}Q�o'�*[��Z,3�ǠQQZ�1�l����ǷG��x�Ɏ�S�c�墩�4�)�k�Fr;�2'�-8���~�VXn+1°���~� �2�|@����OO����Un���n�E�[�&�j�^K0�M��2���a(Q�$�q&�?ш�����H8�ڥ&�A�Y�J�ރ^�0%3V{���eidd��B�B�GP:Z��ؔT嫚��a^]�'��J�����U�׷��<���٪�)/���_'���!�Yq~R�z�JGE�����?t��	'�m2���z�vYG�짻��h c9��Y�;�ǿZ]�RH����x�7Ce����j��Q��yd��i�gGӺ\n8
ɢ��4��f�����*�Rg�X��˒��6�����ި��E�{1��l��j�(��oaۚ��aR�Z���.h}�hT~r�~�8G�b?dP�:����з1&�඾�σXch&��8(��	z #t)��f��4�{��JL�i4���	�����8����#��ß����[��	l�i���r�X㔎;j��1U ���ś��L_]�i��e�j��'����R���P��VUq�� �"-��DѾ��wF�59���%]mܿ�S�6&����]�i ����.;�<��Wy.�ٽi��y`$Y[D	2,���$ڙ�����6N>^�_��5�%}q�,�u��A�>Z��|��I��Sz7�s����hF;�:#7���S��TŐTQ ��V�P�nՅ���E��b�4��V2��6 �\<-��Zo��\*4m�1x佃P�f}4S�����[���r�ןWN�.�q"�`sь+��gs��S��?�I��媺�ɖ<0H&����%(F��|���o�.�O�7�O��l�����>��	u�36`ֳ �:ب�Y�PUh{�/�Wӹ�g�J�@Đ���7���극���t�:��]�K�C��'g�'}�����F�M���M��V�޿]|�U7c�=u'��<� W/xUY�T.��爌��v�H� ;a������^p[���v!���(Z$����V��ܤ�w�@x��/q�
K�):�5�UBBW~QeB�	w)��J��+] ����ƭU�Dz����Y0�?\ͥ�������]��/.L��DU�CNtYj�8M��~�C|-�M+$F���'�ǃ�W��PW2�m��oX�=��oS�,]u�'Z:6a=J毒)'.�]����`�-���V�C���� .d;C#͓�uԋ4�jx�߈����V�'��*4���7�`m�y0�JF�����4�����z2G)�@�-�V���u�c�� ��e	��6����3�"�S��ʱyF�/��k�G��n���݃Kц��ZZ"o �U5!��U�Ŷ�P{ϔ���#z�qN� �i9I�Z�[�R��4�:	��q!x�x����t���ݩ��'QB�>�u�lv��Lʖ*NH�>���ɭm��e\4s�����i�1ᒣ�������V��
�K�
���a��K�Ͻg8�:��E�`t('�k������XFG���cJ�&?�!D��������ef���و�NF�!)�-�+��XlTɜ	��[��N�5�:b���B�O�n����8�oޱԜ��Ц�9���-���y�*j�����t�Y�b�`�_�G���	J��M/__g��gt�S#��"	l=�2���/t]�^f]��Ѥ����bj�f~�)K2��r��3�1@��_�XN���%+~�<�e�&�9�srK��ah������1��P\�ݪ,}���@��a*�4��8���`=T�2��21���,�j�^��"h��S@���a#!�D���� 5��=N桢�f�v��`K?�͔!�����U/{�4'k�le���H���Z��~{�䍘Tf��A���N�pUk���:Uu&~g6ӑ����;��D�ᖶ��o����@�i��W����3�h;~�"wǖ�I�A�kbB�6swv���T`��A蘟�J�_����[ql� 4�: �с 7�yO:q
_�B�ɽ�^��g���@>��{8d�4t$��� :@|�� &�&���&�P�-�j����I��a|���<N�&zۘ"Ǻ��n\�%iLإ c���Ԅ.\޷:��o]�C�v��5BFg0�牴�F��vx��.�+�i���q����tZfT�Ɉ��|�y���lN�,AQ�q�R ��'�>��v7
=<�z�ɀ/�<�y/�8"�/zUB?6 �Ol�Nx��Yɟfb���U} �,�v������ێͩL���Z�q>#�W�F�n��C��VEO����c��a[ȶ���nWN�
`�P��LFı����J���'�C��TO�X@�¿3gnN���Q���!��	{g���y�����wcMz(� ����F#��ڑo��d�
������G݌v�s!��)�:)X�t%��
|d�����ŷ~8�iR+0��H�zI����}o�i:��x}�b\~ƺ�i�Q�����鋐c�nK7��bHDb�9Y��dЙ���ok�8�P0���
��'=�וr��qE�����b�^��}^��7� -�I�r�&V3�>�W,U`fP�� �Y�>��R�z%+����]�"�Ο�2���_c�����>�В�V1�Uֿ�G�鴇G���������{"�u�ٓ�PH�i+����4��͵
~Vî�
��ťV'��R�
����@��#�|{�GDL;��J��q/��.,���SP��k@���W�81;?��!U�)|�O�o���U�����ڷ�X�@��>_�E?W#��|�ה��Wr��ܿ������7/�+5t��=V�O�QFG�~Z�+��D��9�nC6��~�n���f5i�/��͸���G���oS��������{1��)Ч�D������(�vu���B�Ķ��Z��w��ܧ�"�X���d�D��8�}bO�[Z�?)�L�����xXdHx������w26�Jҁ�K')~/F�9���bŮ��2�8�|F�>�n���[*hv���Xp���~�V�^i�d�p� ���+�uWގt���h3PĊ�N+�UZ;�g���\ɧ^y6@�I���.�9����>ДrЋ�� �U�˯O�4V�DE��f,�D�AV5��!B�Ϣ�č�E?�:(�B,��B�p�6�8��ӗx��v��Fz���.���`**}�P8>I��y<�L��W����[�Pߡ[P����96Id���^;[tɭ�CkCU�6A��$Բ���`�X�bt������7[sF �M� �
oz�_G9c��G��JIgNW�ኛژx�)t+�	�Sr�lɒ����6 ����
��T@==
hEs��;̗��h��6?�F�,k��'��(?����Uz7��a���p۲�-�@X9�h���A:?�+�@�HE�;���k�&ɕJ�*lAT�$�L9��F4��}.�wB�Q��5$�qQ�ZB��C�$<ʯ4r��Y�*G@��N��˝��Iyi�c����w�Q\���6�^-��_���!2���U6ې��ѧ���b �±~Uݶ-f ���Y�Ȏ��	E"LO���1���TpK�њ�d���~v6�2��C�3�DTE �I��"�L��r[ۘ�Ue��ɍ=[�R��&����C�"�\��"���'����Ŧ/��v�M��LrPj;{����`?N���9Z�l0צ��fG"p�K�]�p@�n�ʑ@�13��jV�^K}��7�k�����%���0J	���|��3G�3Aπ/kv���3��Rj�ցRA�w_�@�3ܼk���.F, �F���`����"�rEm=f�Og��N޸DB&4���9Ƚ�P"n=�e�{X���'���Bo��������{?m#���-��b�xW�<��T>~4��Ea*,�_)�"@6�h��P���f��f|�����VY�Y�$������ߺp�����f(+���'��TԿ�#2;��1�����88pW�`��5��"�<��A���+�ӛVJ�=X6��Dڣ���r�m���H"�M-K!����W�k����{����&�F@3E����GO<@0F�-�H��D��Ive�7����ӿ�h�#�YT��C�u�Ts�9�ӄ=*�����.�Q�S7&��|�&�V5�����h�U�[�S�Y�ԅ����٘O��}ń�/H���|/�R��H��8�LS��:J��U�B��n$��SE��#��	���F�*��}W!XH��c�/��_�e��@M�BI��'B+���k�Qj�(q8g����R��e�*�&����!�C��b�|���e���e+t��5=GU������|+��Ka��:��R��#��q[NC.T��� ��2��4Z�}dY�1�_��.�����v�e�o�>�E�7���UO!���ي�\��ܾ������+�A���S3K^b��y�fx�L1���-��&zR|�_5��AL�yW��si��3�
�C,�ߵр�	�m�h�&���bx�����g�k|,
\���4UA��RQ�=q�p>��$���h�������+��U����F�Đp��K��<\�������ճe����<�Z�A\i7O³�m���;�໱U���U#��q�x��{��6��e '�����$���_��*]�/j"w4Dr1���89Y�56�]]'��^5�nLqVдR^���3ԕD�u�k� ����Jܪ� D�=�6ER#�%��˩��܄���h���6W^sh��Fqui�ў�FH�J�y�boY�~ZX[��z�����=��é�V!Ă�������t����ha���T����ɝ��vs����AR�r�~ĺT�s]�G��YsaA���kcSB��m����de�׃){V ���`�ze��bK����ɘ�����@��g�0�:�wz�\��-�݂�v�J���y�@ғ�D�w�;wyL�����5���Ziw�(f�&�2�JG](
?3=@�P�=���
,���6��<.��FP��5J��Q�i���H�h�p<�L�=S���Y�s�9W�L�=���Tқ
�����U
�fȌ�f�N�HZ�Q�{B�q��v~]����M�}��ټW��6F`�s�2���[��_��Tڲ�s�Y��f���T���W�B\2�9M"^*�[���.�iB铒3��Ocl�}��B�FW�Z�������6á���G�sx���d�)
XY�k���@�iHS3�k<� ��kK6�t�L�AW�FU�(��GL����*Ag�v�z�)%D0~��UƃGhĔD��4J�L�& �QRC��$0��Bu�v�%N��!��zp�H�ַ�
&�a�ih��P\z̫I9<U�a=�^&���}#�LT�R��hF����x�xj������NГ={��7X+�V��L_t��{♱�n/�]��9�kCb���cSw?���#Οa�N�����on��)� uy����8C��RuoWd�N�1ﱗFH�S.�p��D%���Ϸ��p�3�j׷x�;�(r��C�a�1��MW҂��=g�]S���!�H�Hn�/�L�X���]]���U_�^j�~�%ݓ�9p� yݜXC��0"StP�қ?�}�L̞��TZ����¬)"g'��������]�D3��зJ���+�SM�m*�6prqF��X��G��2�{��� <a���sZ�'��\#�oO�;q{lz��p$�|�""���z	}R�D�ʋ���`Ֆ�o�*�]��Q�Y�s�5ȍ�:F�#�yO$Q��䗟]KZ���l����`2����}�y��ƴζ�%���u��}}_d���v�K�@�ߠ��S6����̲�.�7�4�I������б�3�Dqd?`Cy.�iK�U���a)�iʂdgnĿ��^����,� �8�L�dM���W��!��CD���ǝ8�6���B�{L����s�������qO��ߓD�\Z{���w���[%���ѽ��:0
��gƶ��֩T��#�èy��CH�$fȢ����$��6��6��Jc�j����-A?�\��b#��6���E|�%�����Eb��&���ǩ��O��WV��5����~�)�b��+��j� ��{"B����7��t�n6���ް������΂�z��t�\h��&�S� �\��]�[c��pf�6�Q��Y��j���m�~ْ_jCg�fV,�����@�*8�6��/�s��񶮓�ݙI�N�>�3`��F��۰	��g;�,l랻���3R�I�����������H��8��zԀwE2��վpQ��2��QR"�X(-�w<S9���F�[CW$�I����K�T�<U���p�����bd;F|'�iۓ~'I^�C0��u�ǺgйmF
1u�/�4�4e>e`"�TN�ft�`ЊV�B7�(��U7�h3�:�
h�zdx8�,+o��`X�
�zi�0�~�#���Z��G�!�r��Q_�\�5�����z��p�)��x�c)�s�U�/	��嗼���F���������~�O�T?yP}��Ycq� ���An��J���7KQ*'��+viM<	����`رc~	./�ݡE�s��z7��ɩ.�uPW�5$+��&Fj���T%�J�kg�P��漰�Q�f��k^=�&�To����}j�C�Y��^�|�8.+5F�3a����Xg�<H���[;�:P�Ѧ������a ��[�/�<��y��G��S !��ǂ��?�u��#���?yZ'���B�6d�&5��+�z{�$B�ZLPQ���M���$4�AvJ��Y�c՗��;J~�J��j4¨��di�Y
6�u���X{6]>���Zy�ljjS��w��Y��>�Jj#]�)��o���}��-��-l�ߙ��n`�7���}mR����,:5�����w5[�����֓��[Bp֬r��ni�Z�����Y���_���_��=�A�U&#ӂ���ko:����ԉ�ωh�g�o�x/>�h����m̀��Y�� r�蕶�'i����F8�X�?����s+Xz��k��fS6X�ٙU�������昝C�/k�hD�U2�����w�f� �J�"v��,D|��t^ �͞B����fO:L�� �{�57���C|�1��z[d�q�	j���xI �7q�4Ns0��13�f�B�^U���;�>ҰX$H�$���ʈ��Ym�!z�MӢ��Z_A��y,(u�;���bܑ7�J�\�W]A�Ҋ� �L��{�D7�Kn�遄O��gm��2� 2 ��$H-�J�e��G%�"�*�ና����<Ǚz�G���sm��y�>^��.
n�g�~�����
��*�}�-O䈯=k@2~0���x��46��ޛ�NW5���u���i68�"��~��QT�I��q�[��I?h��l.6A�o����J7�����o{�u��U3ꊭ!�@�"Qh'`���ۜ<<����EX�v ���uy�lM))ǝq��dCG�ZJ&��ѻ8ժ����$��Ua��vM)�ѭ��n�-�;VZ���t�3�h�|d�+6.����-���+�t?R"H%��)i)�aU���I�F��7�^"����������a�{5�ȴ=,%���6��c[������_{a;��d-�E�vDT���{�OP�|0G�W��WYH���l�K�3��4j���Ne��3gN�a�>Ȑ�X�&Ѽ39q5��/1G���a�����Fv3KH~�Ϩ��&��ey����^	_N��6	�V�<:M]s��q�"�;T�_����{�:��'�Q��jeV��5V�$*�{V�{>�;:@�,�VbfA�{�.M��~O����S2V��/i�_��8��iU�:��*�ۆ���
4%R�D�@��u]���ܢ }����𔫽	���E�Ϻt:����5�kfE�^�Q�%�����Ә� ���z*S"J�T_:L�O})�]�ٛu[b������X��`����^r�Qu��ǹ�^At����e@�c�H�*�'�|t�X��y#^�3�y����H�����]�1����c�r`��
a�>����y����K�5��m//��u�R20s��ݩ4S��BO����[o����8Z����v�\�_� �ve��lP[�̣�c��D�[�u��Q3�c9�H��QطM/���Y��d��Ն0�C�����3.u�|ALQ�ن��at\���m�ӻW��o_�i5臞l���k�io��)�͌&ՠrt�j���#DJ{1����� }u-О��O����f`�f�IoȮ�6��E*Xpp����=�L5tE��V)*���cΝ qE|Դ��N%��J�K"�w"���q�Te�d�ːnG��x��
