��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����0� ����遼�6������"���#�{A���'j�Qj} �}xT	g��F����a��f��洜K%g==�Z���L1������bG����XB�k6T��w+F��3r1#�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>c��mW���rJ(���/	���~J`2F�x���4W�0V�y��l]��X���8D�G$�ۻ��c��rk�E8o��W��z�����O�Q�F��?-_�䰹��Ny����o��:���l�,�:^�G���G��ta�`����k�Nx�YfU���}*���9���e7t�T��Y.�����y�0O�g8��B� '��xJ�`��M�w��B�H*�y��MkO.~�u��6�-���#�w��M�#�j��!~�����h��qf����i��&���T	0nL��J��Х�w�r�2`P�=�"O���dB:�&�C'��=����'���M����wr��i�	���`��S��s]�_ה�uh��"��ܜq�0\���t��ڃ���r��1+���?�m�8�n���Qh�T��Ep�V�����Vo,�P?7(mb��8{>�"��Iw���D��NI�G�M�!!���3��N�����u5kT>ٻg����}6��PUT��y����;�9p�<�}���~/o��]d5����p�/S�{���b��w~��1ѡ�,���%�!��Jbf�\�C�FU^ae@��н����-�5�f�Put��J�T�If��sޤsK������]v�+HX������p�N=��E�rҬ������~'�=�2:<;�C8W�4n"�n�i��q*o��]D�A�]iַ|�
JI'K [�M�{��yRO�p0I����y_��奮���ֹ��}I��%�B
	��"�^���}|����Լ��x��j����l�E�{���P�e����.��
64�Î�~�Pb��^y9X�N�g��� ���x�O��݁\�G"�B2�k!�i�N<�����2ɳ�\�n���ۤ�)�a��	�8���@E��o�����E��*B��Ѐó^Y찵̸5��ң�I�������RX�N���r��_�'��B�\�����O��/\ʘ�6K�W������C�f���e�NS5ʧu�'��{��*��@ A�W����vi��U:���c����}[�j�@T̶R.Ž6�������X�eo7��g[����(8�fZ�Ų�	��/\Rm)�JOS�fn<�t"5s5ƚ� ~LFg�.kw?�К?̢��h6�Kbg��d��#KK f�����(lNX2����)4_(�����C��30�{EM(m�(�Hx<c�,r���g��Q��._�߭�0�T�ifH�/K� E	C�s��?H��iBkQʘ<�s��g�8C!oļ�3#�y�����&�[�J�8�}L���ڦM���3>�&ם6�"DHa#q ��{*�Lqe/����K���qS�e��)2��M����a+ز���c�Ri���GIFd#����D$.�c��r���s!^�������c|���_k�|�s���l��O��u���%Q�s�+1��8�(ŵ�7��%����2?����_m���:fM��A鵗�&�v9�(��]�-�G�{�HP�zqg˵����V�J  !��Ar���?T\8���r�l-?mh��A.�|�r�̩��s��8�9�я7+ �-�r��2ϥ���i���D����S�'^���D WC�� ds$��c�x��'���n� M��JU���Mi!����e��� ��&�i�P.v�a�s�Қ���<�*��.���dO9W��t�1�I~^��/�'߇���K��I�Sn�G�BBӣ��r���Ԁr=䩆�*�U�t/ n�K��Q���{[������n�xY^"=l�=�-d��^�a�:6H�G;6	iqtryҙ>ŵN�խ2}�@c\�'�5<����	���X���0�w�����>��v�[��,ʝ/��kw���D=\~�.���4�K���V4�W��WK��fBм�v̗e���I;�U���%��2OKL� rPN&n60��� �^�NE�kH2X���g�z4D�Z�FyL�n�v�RF2Ma���
���5�kYW��7f�ݟ�����҇\L��>H���B�9~��ھ��ZŪ��1w˰�}���]�]G�!g0�[7�a��	��T �"=����Fh����S#my�EL�c�>��j�J
�TO@�(#�[W|rt� ;��ĉ�I�[��4����ڑSқ�qel _!bƬ9z�I`>0|@��l��]��yZY�T����/==a'붑 ��-��Q�]����/1�r�}����3n�л��`|���x0�A��j�*�z�p]� Ep�)���F����o2��9*D�O1�u1��ԊS�;�;lԧ�C�����w���S�� tWEn�6�y�-����a�o=AҀ�E��&;ʘ���kB4��0f�v+�?� ��� �0����ĝc��>Ͳqo�9lʨ]��=�I�Cy�M�dHwQ��JI ���d���Ǘ5X�ڜ�pl�{@i6	���M�?p�V�]�u���;���L���wS/4*�8� /ۀ1+���ª�R7��:]༬��s�Dɔ�*�ez��$L[i.�_� �d (�K������Q�%u��`�4<N���[	66Q����u�����fW%�_��/��t��E�۵7ZZ�k��X�Tf۟�4�;�$A�ga��*�xy�X�r���d����"$���ą:
�~�ݚR�K��v�Ap".������>4�+��t�h��_e�WK.����{�D�ؾ����$!�ru��t��\u)G�s�?��^�<j8?q[ku�I��-� ���|$���pVg�ߙ���"73��]_А^r����53�K��2���ʘ~��n�	م:Hۤ�f,�
���;~�� 9���� �⍹��}��!i��58K�q�}��Ir�z։O���#�����?�L?���E1˄�/��\����A�q`�w�_8���1Tџ�)K�'T4U���������Ny�E�~�\�������8=P:��l�@� ��G� g%އNR�q�
�8���l�f��.�FNK���A���>��ž3�!���nXJu�t �vn���iX�X�Vi���~	�;+����k��OِL������z�������%�3� ��ܶ�X���i�J4�W�NT�W��t��k,ݩ(�1�ȧ�1lU^���B/:�Ƭ�O�*���)���ވΨ9{
!�0&�b�5a�жR#,@�s�Cd�)�X6H؀'7�6y�_���b��d��/�-�t�G0)�ۙ���JY ��]%�Yﴐa��Tl�G�����:��a��M���� �j��r�t�,�Wшi��}w�Jӹ$Q�4e����> Fdv`�