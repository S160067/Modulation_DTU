��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����0� ����遼�6������"���#�{A���'j�Qj} �}xT	g��F����a��f��洜K%g==�Z���L1������bG����XB�k6T��w+F��3r1#�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htdʮz_�0�`��@�[D˂8��k�ľF�n�Ԥ��r�τ�u�&&����\l&�$������<H�����}�ƌRS>�(B-~�� ��ڣ�9#M��c��&��C:��p�@n��7E�wJ�h�F�p7k�=f`ez��1���d��D9��*`������t���篞�JM���8i�):�ͦ���H:|>����!z�ml[�<�a���Q-�L аz�H���QQ_6�Wr�,O]��S����~�ڳGyOFgOzf�1/�]���k���
"�
��;f7�/�e�̟�����`�E
f��z�m��R�r���w��kU���KV�ͩw��:�\75���E��ڗ�p�[�u~��{E�!�P�fU��/�l�<E����V��y��:�hA�1�����,�N06�-&���ȴ���F�t�`�X��l�*�xE'e,$������ ��7��=�j���A<�%h���]�to&0�� ���&nF�O�r|�����>�����#�1tD�k�V����N�@��n�V�,�?��c�M,��	�[-�Tb7�o3�&��戱��'�T-{���Dusp�o�����Z�:����������S$�p�
ӍϘu"���ɧo/H;'���HĴ9y�'j֜�I���z�Ws��q�������I�.o�׊Aо�vр_B)�d��ܸ���=�QH�ӄ��@���(kY]�~����M�������n͹����	e(Wsx��̣��1%�$��M�Y�4����<ӄl�W!�CP���HQM㙋Ͱa$�ƨ�b!9rh��$KF��f��}:�$]�>(o��I,���vD(�w{�)�1��J4��^��,��'��f��t.�����5ݸ�D���&�X�4��X��9�@:vR�ր0-4 n.��M.�����d�)6��tT�cw���F7�����کή.�����$��+�L��+�i���������Vf���:���;�ܣ��u>^!
��Pv%��l�����vD����/��Л�\9���fjMo�a�sA7+��#sZ@�"�W���� ��'��٨���V�SG�Y�9Z�u_�1ÿޓ��� H?�q$�(=�K
��BF+�A�8^ɻLQ��6����_������)�6,/�y�Z���si	߈�����Q��`HWv(ٓňҡ��(?f�*�I?[��ɋ�*0ph�D��by�!�g�r���hX@��n.N��>]1ռ��U��t-ٯ���(����P^��}D�W>Yo+eg�o��w����T��`
j{����/}3��l(�X��{����E.�?|�D�/�GK�j�-��}��,����� *=��l��
Ub������'��kO!��V���A�ِ>I�]mRB�5g��o	�� r����t!�����`DF���O��_�$�q�C$=���I(D�����qm�NG]��=U�Z]��Y���AW;�g�Z�������?E�O��BvA�����[��s���:�k��|���/h�N����G�� �ˆ�)	���V��eӛ�(���#6� ��Wk�X�Y�/q1y�7 a���qe�?�|O�\;h0��O,IZ&���^��F�D��/~�k�CC����*�,�.a�u:�cŴL$�2Ne!���ٲ�a�~=��#uJ���)�f��6��%��F8�phD�,F��!4��/��TY^�	���:-�^#�s��ѳ\�8�A�C~�J�� �o7Dhb$��h�L�.�i�T�!8¯u��'�o[��ՠS�*3�2��d�E�W���P��j<�FA�	��Q��no�JE4z ���n���R@�j�K�jun�	|���Հ��z�S�(�)�a���������Bf^m���:�l}.?�y����w�<\~��ǥ�hbD��w��e�Tm�.v����ߺQ�S� v���״�~��i��3a�H9�H!qs��jo ��"�w��V7�"�l]�_��W���A�b�u(����^׎|'�	rq�f�w��1��?u-2+Z��+�T��;[5{S �h��i���ۿU ��}���Q����<�Y!�s�����O�e}Wx�El8���-�z� �YustM�-��rL��{�*X�y�W`��]���q��~�V,�v���D�^��X��r^��:�*�:����7��]���AƎ�#�O�G.ń�O����R���N���`f�ڣb���<	ԧ���bik^N���
��<��C�sq�=��IϦ�).A�b�����~z���Fxez��|o��C�f�JNG�� 8W��0@t�D��ē1%#���5���3Yvc��q�/g VΔ��DP>��z��Ye�/��9s��������'�6v́�N6f�d�0%B]u�*1����0ޘ_Ig���T�I�j4�ړA�Nn�n���N���7F0qh��{\���)���D�j��fVL V�A��|�ei=;K1��Z�m���Ǌ@>y@BD|�C���%��q(��f |�s.j���L��[:nO�ِ����Lh�uabtnN�����9]�����9V��
�.�d[r�9���[���ؕ27%���I��>&�������&�]����?;�I�F�I�
r��Ӵ�=���G�&��dx�ux����� �P傗�gx 9��ҷt�\B.�>��I��H!�G�~� �G�X[S�p�R�݆|O��T�����\ Wv�a.n���J�4�op=0N�(`&F�+��wd�&o8�cɞ�S�\a9�А<-�qh28��sX�2�
c��G�o	,l�N���?-����TC&��d�T�:��5vd<�ڊ3�Q�(����k7�Լ�G��O֥?��R�E��N?n�E����B%tsGE5��|�x7�5wT1�s\�kz٪=#��+�('	V��H������h!l���&kq�3^-Z�f�EӬ(wr�!�����UnU��
��s�+e_)�h+-�+S��&���B�H �77�����2O��l�+J������hDO�\����?˚}0Wk�e�T:�}k�Рao&���j�Z�b:Q�pr�BEsJ���Y���C��X&t�8�ȣ
^k0�G�.)����a;B�/Th%�b5��zN>�o�H�x�c�ډ;-�e=���Ѷ�P��,��[~ ���Ү�t�V�|��Xl��#敻w[2��'hh���i�y�{��Tv9U�x֍?I/'� �~����R������