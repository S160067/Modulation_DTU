��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����>�S��fI#�l7x%���$or�#�6�y���N�i� �D��f(�:eǊ�` ��S���^�mBƱYjA���v�0��kh������#�v�(#W��ux��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�O�AC�Dl�w��;�|�y:�	��gL�0���\X��D�0c�8�p��!Z
�O�.s�H��/�hȍ�`���@UR- �BϤ�YgP�C���/7|��
���EM����\�Ұʝ@g����JDyܳ�b���bH�7a�ȳB*��S�!0�PDk�|�U�S��D:�Gl�p��q��لe㷗"�Cfe��b�ߺᏻ\5�2wϺĒ��S�;~��ж�Uwr�ޫ	,S�'>�q�Q�T˞+�A'^Baf�AC�1��~*��W23�B!�->n��$�-;�])x�Qḡ#ۂv�֌��䱥��o��n�^�_YzG�1' h6���Z{L~&��<���E���h��Ә�7���&��qKܖAK�����] �� &͢$m`�&[(7d��2ȁ.�i��h�Μ�r��n�2Q�*��W7{��{��-�	VT�׹m�א@�e��H�;1uW8�|�X�"�l�[�����$�c�@���-Q�}񆖕�k78���^@���F��B4�q�(�o��� �!���,@-r������Fa#L��dO����`.v�ћ�2��s��*�Ћ����9�-]+}8=��
4"�8P��<�1"t/Hxץ�}a��`�ª�&�y܇f~��z���Hԡ6���Њ�1��K���/�Ң����Y��@$�����T�*�x��^��jܐ�$������=�U� #�(�oS��?�������ڑ[i(q �.Ai�o���.�ܜ��n�@�]�+�i���+D���TU�ܰa��;=O��+U�h����&5K���������K+FQ� N�T~ϭ�Rj�_J�zfjm��X�����}�����i��!E{1-ߟ�t4�0����JJ�Y�۫�2"��]��q�b�lZ�w�q�lF .�[���H��ZFr�=�p{���k�	�7�� ��%B��'�ȝSGff�Ta
�Z��8+3+ʃ����>3���>S�� ���0�������
���u\��P�%��=�1��J�A�C��}�Z����(�{�'|�� ���:�ꂝ]s�c�:�6���A,4m�	tD�y�GOO�h��w����t�����#�	�?�a>����q�~'�*H3'���pK�Q�*����b��a�-޵jQ�|��4�|� �e�*�NY8á����5�l1j�	G�����;y��D�i���-��i�d�yx�v�+���a��}] ��	�~!�i��=3�*C��n� "w�jWtPs}E���T֛Y�ּq�eͫw�ӕ��R�U��8o\�\LL.;iO�#z�8"2<F����=�A4#i`\��j�
`�Y�K0?�W��i�����=��$�c�,����^a����`T��= �E\]1�ΉN,�}�K��]�Ǵ�'o��-�s7�%� M�m�%qp[���%E��PK(��Jw�*D���T�0���.����5�슃X8��'~�v������=���Άw�n���	gm9�S��.(8�,hD8�B4a�S��|U��X{oS�����Ǘ1��-��Y���������H�í�KyR
��r@��ҕ]>���.��~������V	�o=���3݄��T�!��h��M�h��9Rd����3P���s]��{pO��eѽ��+��et���3��x��o����5�ɐ��?�]�?&Xe+�)��j�tg8��`��h�хs�EfE�}L���{lD&^�z�q�C����<'�)?:�a�i60��sq7*F�n��r'-<������
U��jֺk�}��z'�=��h�H�_j�LZL��S�m6�Eɴ4���H�[�ϖ^�K�~�rg��<[�_A�^��	��h˘H�-��I#\�B��"<��e�y|�tW+�$<�@˂f��5�g3�l�zV[����1+�xp����a>d��ʐ�L�Y«�~�����>���΂#:T?������������"��NN
z�Kb�:"Ѿ�������� v����C,�R:oL�4o&�� ?ܚB���Ut^I��f��mh"k�f3p7{���9�@2��#BѾ�y�HL|�R�*^�"S+"U
Rt�,����ruq��hx�W.(�5x�/���^��Q�Mad@N�����o�j�[ɲVԲW(Z
���0j;��\ݑ���e``Ex��P�nqE1�¦�  ��D$6ⵣy��T�
h,��S['zu���(�<�`J��ӏ��"��Ea��=�N���A ��� ƣe�����i�4۟ݴ���N��.\���#5�^���x��)�����X�e-[q���G�fү��T��L�K�z��������\Ti���"�HdF�c���~�xU���@�F]��/h�> ��y4O��"ZӖ5ǝ�+dm��-A��ڒ���H��X�0 �^V)�p�Q +S�+]w��՘(w0�jE3����&"���d�(�"\����D��7��4m�G"��b�\�qM���"2�� �>~����_U��߉�&wN6`F!­/@ʲ�A.�'�ˤ���Z�M_/�]Z�6z,�B�\se���2$��)ʔ�`�͈��|L�5�WLb �h<��
���'!|2��>������6�T1S�j��7��N M��9+ȅA�T�n�PWu6d��h�=V�F���{�X�z�=!�8�|���aE҈�( 9"�Z�?�c�_���� u8��'0��cm`B�NEn�J;���28�����7e�Y��-�V&��-@_qt�P�j,�p�/z�,��8�Ro��
����֗]$yȆUX�<�d��s�>�Z���v߾-�[�(ߗ\�
�:u�����Joā���9�*�h�L��3��˕WEp���7?�J��x�:h�Ζ�S��U�LD�?~P����-[�,�ՠ�J/Yin�����a,k���_�@���1�����Y��:��9dE�!�L!3CK`��K�] q��c� ��-�rw�J��=j��ųȦBֵ�뛑5�}ڰ��k�+v)�2 ���LX�����g�n��IP�r�%��ߎ�|#�{�E,|kw(LM�P5����Y��<���İu�Tjen��RR!�1�@�oΟ�f�`9Qvn�$�΍��s�v��P"�zwW����f�h6,����Q������ce�kc��٣��Vˊ)�؂�߃{�63_u\��KZ|e9���U� � \�8��~)H�0���Qh����D��tm>�җ�YK���`"��3�7���>�� �gvV"�g�����8;�<歵���5���:\��/��'E�Rfl�In�|����w�5
��N��W�5˦�K��<��'A�Y�ӫC-�h�;�;����(�|B)�@�~��?�
Y� z������T����&�8�Cx��az>^;_�C�-%
y5�����E��*������͸������5IMA2��f\��@��G}�["l�O-�w������8�-oa֦��#�f�:��'�i�E��c��JS_34<C�@�wȈ�e١<�;s�h����`Kٚ��;��ʱ�/W�Q��bM�*D:b�P'k��*�
����$,pW(���=Ӝ��+2�yɭ�_tiu�~'��w��:3_���Ǻ(X�[����|z�5٧�)D��o��P��`!Y�uxP�2�p�����h%6�5Sͭ��尡~w��}��Y��7�X蘅���.�W_d2��)u�L�[1�q��EH�ʦ.+ O'����<>l�!��
���|=.͝�9o@���R�d�LD����?�$FE�z�}�~�X�p�����@f=zvD����A4���"O`_��n�+`
�����@s�y�n��d�F��(�F�R"�q�`�"pd+�[�>.�AF:�sk����S�}� ��'���	.+-#w�NxiC�'��ZTb\�Լ~�❾*�o�H@��`r���|�L �zӭw�k��8B�?��¥=��C��n5l�ê�m+��~T�s�~D����Ƙ�L]�*�����E�|�|nN�>$1���epʃ�W�����	[��dPTC�+e�*�ƒ��p��#bqKZ�3�S��VǕ�*��ikH�s��G�������+�\���������,�Mos=GE�z�3�X;�1��cd\"�e��ꛇr�#}����
N򇃖@����O��z�-\%Jlg�X�ſ)|L�0r�zk 6�Ww�<%!�n�SK�_��믠�\�@�*T�u|Q�T�����Z��Ŋ*u����y�����}�P2Q��%V~�>���%J�ryt*���4�]�YS��z�I����s��PJZ�o���sI��ZnP�_.=�sMb��W�A~�S�A�X	�̩$D�>�#���^�Ө���|�ܶ�䅝�P�-�����F]^76X�+A�$�o.{F���S�ٔE�aV�
���Kn�ܾ�W�J=��9q$�3,sl��Բ��I��ߔ��ee�?��9
��j���J�q>� �HeA@i��鑵~f�
�B�# ��I�E��,A���B*�I��7k��U��|�ƌ 	\�i|��y�E:�~x���5�+H;d9�1�'��O�K��*�y�#�6B��B�f�u����pQ1��d#7��%F�QL��V�t�]]��$�NK-�1=U���KS�0}¡����ֆ���3%li;�@ɍp�� ��8�ǼŹ)\�AxԼ���lA��"Yyww[�R�c� Z����X�����HE�F6�I>/�`�@3�)c�2Z
0���?@�'��X��:��5i�)̦�+ͤ���Xw��.?٪�Q�T��~�����_Q-�%8ǻ�� ڑ#��)�t�m�C"�x����S�L��"��� �ѴB湸T���A��O#)�,O�c�c7�ځt��S�եWh�i?��q2�Ҹpw�����7��Y��í(���7Ӆe���7@����if��k��j��:�3��U\��<-��6XUY�rN���f�L���v$�dt�?�-2?�XU�9��Th0ɀ�C�y�p���e����L,�A��)��.�/��q$�b�a}/�ނv��E�9l�w%��v�J��Ն�~'x>�5���z?�B-�<A�)k�I�ӃF�}�4�O|E�(���􋗴t�������K�`K�,�Ր蟜����Rf���:�}�Q�8���o�cG,Ey2�U�Z}�󡆡8A��#�i��`ԪʜRGL����dp�a#?��ɢ�X*���C�.������NA�:���<��a褮k�}4��τ�@5�2�5S�Em���dk�eJ��=d�L�3&J��Ӂ�,-@�=��rs?Y-�U��S��Y�q�&p���Yh����q�_��0'7�9��?���y;�Jj�ށ��U G�3m�%{k3�,��V%`���LM����z=������:~+�?�6�\9 �L�:��5��8O �&�Y�d��O����}-��ANƂ�A�0�7�m�e�D<T��=�=���?n[��il>%vΞ�:�'�YPA�t���K��7)�x��R��:����3�EE%�~�<A�<���Y�k� Q�$+Ɏ��aS���ŧvcD~N�.t�R�@�A̜`T�7S�	���*4I�4N���N�HQm%��
W��ݤ��a#�v��0�ߏ�u��)�~!�C�yD�އ�|�w�$�	f��M y@
���ے��U�ީ?�B%�ٰ{�G�<�<ā'�����<@lL��hB�n}�:�!N>w�_��p�<6 l	M_�^�[�ڴg��+�ta������׺��9㨸���j�T�[����S�����s9gp��sfe���@,��?H�4o�6���S��8K�i�0��}+�N��/Ť�Bw
G�,����#��8���M��� )���8���|>�\� �0~%��EM�Κ�??���Y�� fS���y��58�� &�.��R�Nx׀�b�$Ք;�t�B '��I=����Ʀ���/ ;��%�8��>&!���)p����+���Jr!
�2;�b����E,{h�I��s*�a8��:[Z|+��S� ޷������;<��d-XS
^ո�!jb���F��'Q,,�*QA�r�	n�T(귩I�M	�D�G��Q��h�f��F>��#}�/��R� 7�0ӂ��v[���i}Jƕ�m�x�ک����>��A�@����H?Y�^�2c;�;�8#۝�4�?�p�(Fh�f@�!q�^�#��J���@�yNJC\��(i���M��b��� ���D��)y뭀t~�&d�dB�l=Hb�hC��-eQ��WXh����x4�Dڟ��L�~�
B�	�P�{�T�]Q�r+�^����D�Eb�/X}V��R��GG���;���k��� L,��5��ýץ�5O�<�z��m�;,�u�s�y����c��sW�Q% �gѵ�&��r!a�)�T?t�	f�Tb��>����_"�y-���dڃ�DH0���}�?[L�r��
��m��U�{�
X=��/)e�H�zTK����bNձ�2Z��5��B�ٌ�A��=7!��F$���O��й{�����d|i%��`	*;��G&]��Np�l`ô�N9x���goI@S��Lщ�YUz,�eh����ku����PJ����U��rE���������]A!�b�H���x�x뜅�������)�Ch�Cc�� ���+�+	�l��4/!��H��`˲��������t��H��m v9�.'[s#�0������v(r�Lƪ�4�ԙW�U��Q�%�v�]��Y����u~����R�x+�/-2&4̦�4G��1	�^�k���΂���s��� �Nn9����C}9*���3߯E��1��t�u�!�)gq!ġ�4�_�Q�tH�w���w"��T]�6��$�"�KH��'�0Ą�-��ρ�f���r5ӕ�d�7���V���K��(���ە\[{fwu�5�	�����1A"<���	��x�����!�Ar�/�<�(�����0�b��I��5U�t��+��U�y�^⾙�93�ٝ�mL��8���9�D��4�RJ�����j1؄��.zi���HΉ�s݄50@o�)�ܵ$ ��Q �E��4�_t�Qv���� U�Q�����>54�l��D4�8C�) R�ҡK?�cD1�	�����