��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���,���`�Q �����6�͍	),�6�md|_��n�x�"u������K �5owJh�E��qڑI9����%,%UEwf�x����;.�9��p3��,/�֤����"��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�Oo�Ne�<��!G�u�uO]�nG����W��1L���a�KzܸƠC[#f�0�����-V_� 8T^(�|��Z0��+����[VT`�c��A�p�����	�S��60�W���)/��L��A�g87V�c�5�_Җ��sd�����PA��C%#!^��M[��[C�r��O�k�#H�w�c���T��7rC��i ��)�sI?�V�K7ۉ0���F4rg���W��:����J����Em��]������ \do<<(���1�'��*��{�"�%4P�D��V"R��G�xVxV����\��T:r/����q�B3�z��2z��un/D��QG%�=oTK�;�I%�ǿ���α��|��mی���o������?��H��t�x��M���ug"A��w� ��fS��������`���?��X���N�����^T(�u��p������l�YA?����L��bI���7lc�f�6FnEq��Fl��� ��g�Y�)RyX蚞�u����^�vTC��n���S���]���TWq�x�B��˽{��`��*����h*CN@�-�C>�_i���8_DyS�b�ʥ�^vo�0w�����a�?�1n� ��Ǭ� AR�ϓ\6��bu�_"[�P8p���	��1� �өVt� .m3�p���Qr�%���Z�^��'VHDb
v4�;/��u�_��e�T�ÙRj��]���u]/GR�r�ۣ|w{拈�?��x�N-�,����=����B�H
�b^"�׉��i���+$}\T~YַD�K�1B��q����u�(Rc{3=����ng�8Z���5� ṘB��h��T<�;92��W���}������F�b�I�:y><��#�c���Vn4�{Ʀ1��Qx�b*�G	� ��5_�����քl��l4���e�Iݞ>�#6A���ؼ=�gi��6	���D�8�/Y�ėגZu'���^��YD 0�^��q�<�l�Ϻ��+z���L#�ʦ�LA���d���t�.�PT4"�̣�H!J�5G���zR��h�x���2�E:�X������Ѻth7�]\r��cqc�\����.o��g��J�}"��������s�IY��*
Y��x�v�_�m!�r�֦*TV�=����F���a�p_�	s�a'����z�;��Q��̓c���W���_��L4�ٰ��6�I��GLκ�k>VW��O�Z8�L�d��\Ȋ�l�fj��l���	:��I���aX�`Im����~a�M`Sfp����o��+bCVl0�B2�}�xd��h�EK;-�������M��H�'�7�Q�iO�#�r�,���;A�6�Z���4C?�*N�b�8�bh���T7��F�]p�ȍ���&!�V��{6��%�5�ocنZ ߫���	���Y����6���h����c}�1}A5/1g���3��ݮ3;��lb`�51~ߖ��P��#�N mO��������N�S��8#���}o��q�V����~�u����2���M葊��%ƣbڡ\������MĨ�(�M	���t��Zą��V�{˔��o����p�����F����ƄИ�w��Λ:�A���CR�$G��qK��@2��/����>�XqڹH�X���#U���@�7��=:����D�(�����đ���DS)s:Z�G�)Fa��Y��{��e�A����d�к�,��>
��=���.��L?_�O+�*Y���&�e,�A�cYF�Hm��������͍}hf���YO�����m�߉���Ld��kZ��όKx�=C(����m��+2r�ÙS��Dk`%,*#(����_�;U>���Cv#�I���T�(�y��6��+��G���gi.I��~�E۬�����CS�m=fS:�Ql�<:�����_���Bs�t�����g���6��!��uð��#h#A�}#���	����ܡ�LK���(8�����6�' %�:���y/@�x�`�90�,����Gd�=�g���Ng�JmQ��LcPG��]:y�4�9�DɈ(c�csE�е��sm�y*�˒��t�e	\���;��^�����|��c���n�g��!��&F)3�d��>�hs}J�_+�72|�_��ּ�η��r�3U�[90Ԫ'X�N��b`��Е>z�}l����@v�%����<ֺ�fQ�vl}���Q2g%������z��F�[U�@�j��M:w�B'	T�N`��9�Xj�-2��Q77A��g�Z�i���o>��=�|�:�c ���ﻈT�|S�r�8���d̡�lp��(�wkR�b5ι3w� �U�a]��8ENBW��;�K��9cP��<���[�Ϧ6�G�f�+�J�ͥr�&�ܛ�j�CEa�[F�;īHR)ꑊ����"ċ��!)���h>�Ͳ�c3=�U�>��5%�빱�J��=��*�]O @�pҝe]���ltV����$A	�a��^�K��x,O^������<�*h��h����2M��)lD>�:����Hakpp�r4@��/|��g�W�T�"$�Д��^;��� ��D:�������WL?���LD>K{Y�.�3�I�0�ٝIM��uƘxǀ�t�<Ip�������/�wRo��K��G��9�ݲɸ���}j�G����}�pS}�3"�f���(�SB,����9��[D�K)J�mө�R/|]:T��E�a�(��R�w��jP�g�=K��	���2��ڸ����Nȴmo�'�v𚌿��/�_5�~?����G+Yb������*f�D�񙕳�1�k�R����6�'Q8�[���9��/��M��Y5`��zv���=,�`��
~̭�����S�8,�b>N������Ծ�NnҬ��-P����_����]$Y�>�]�dF��=�d���u�:��tl�f��u��ٓ�W�*/ז���ɉ����K���;�aJE�P��>�g���]�:n̢�}�Y����Pz�������As������Q�y@��\�af�+jR���]�h�gp/���+g{�L{����1�Ѣ���Gg7�����p���XFM����Z�bDq�ڛE���54r|b����?⇦�B.Cm+tȬ��G���+�f�Q=�j�*VZ�����P�(��ܗ0� Q��%�=��k�sD�x�_����=3�N�������.1����$I����@Ǟ2&k%�vm
[�J�����%�gb����;4_�|>%L��<Z��o�(k��l~�߭������͵ߏ'�7����"B�h��鵀Eq�I�kؼڈ!�H����J�+�[A@��%�!�1�o�].��v�TMN"P[��]U%S�0��4!�~*P8��"�]���+���R�V۲�x�0Z��\iS��\�����7j$��S�P�z��f�_!b7�S�ڴ�K`��o�+m�����u�&eRƕ�=��`MHa��w�5�1�X�V����cq��3�r��.�br�rJ�=W�}/!%��O�lߑ�g�ybۯ8)ȉ���<��1���#�ټ�O����S5�t��>�,��C�5�@�7S��U�w�I=F(w�
���a�f���H2.�Ƌ��ݐS?˂d��it;�Q�v��n������,p������d����!�sx"�/UeQ�]�`~�%���7�a�S,��_߄t������&����7F�x,���<%*Z2nT2���m�竗��Df�d���n�[���|g��p�.������T��&�˿bO�tz'��	
���gWǳV��T�����&���[�PI^�P^�+�l��iu`�����T�x�{�����k=T������"�e�%��4P�J� ����x+Q�+�G�\���ʑ*��ɳ��$�!�E��*�ݜ�'���[*��ɇx�Q��?2~�Ke3K�`�/��[L��w7��٤NՈ�p��k6j��/����U�N�y�
,��;�,�Y*oce���M��A{� \A�x@�l��Ңޥ�7M�DW�䷦�>��B����Gԏ�ڭr8 ��h�t���7"U�~��y�sQ����ѿ0�c�F�R���
�A�ZY�Kh��|����s�b�9ꄟ�Cp%�M@��=�����r��FO٧��v��x�^0�b�{[�z,'��w#�ې�G�\����j0��7��>�s�� �y(��qV��O[@���ܒUU��(H�G��}��IGD��C��A�,���*�gRg��u����G���hg�
98�YӅ��0��_�#�#^d��w�Lo6�@Pۮ�E]�(�)'gm�XJ732m�0������f��׵W���{�A_�[�JP	w���2����� T)���K��~k��~x8Ѿ��HzR��s�83�Eu�md�M����o~X��w�?�? �K���� ��H�ޓ�!�ٜ�\��!�o�.]�u�(��A�"�g>=��<6����mC��?QR7/��Gg�,�}���KD�قOb͌qpU����k-���u=���q@�%���xf�V�^�w�`R��\h�>G@�!�n�������x�݈���'�0�wڲD~��ʠ�k����u����1j囻~`��T� ���9��U�E��Sf��P�Tk�I3���o
���qn�~�y�`���j"j�Ӏ`
�H�B���=���8|}%w.�� ���[�h���	Nr�����:@�b/��KÉ�TM5Ag<s���n�m��tz�.$�x?��e�D�u�p��5/�¼
�Z��
�yucPؠ���*��	;���wZ �B�R�H���X��7�)�r�,Z(��ktO�&���<��UL�Üw��iZtg����/1�E�'2B6I���|�2u��|X��ǝr�ͷ�[f���OƧ��i�-˷F�2 9��5�B͞s&{���/�R8��w$���Gڨ�� ����|����:F�3>ڵ�6�']�G��YяH�w���l��f���]^PZ|��X+��X{�y-q��MB�+��߭6wT,�k跤]��u����a�
��D�x�J�~�����SX������{[V!R(��̹�82"3��i�<Å>�)�=B�z$7�-Vt5K�4����žl��^KS���"�ug;�A.��'��F�vD��2�q��Z�}��Bʁ[Z���?�w$1���r��7��m��\?�����%%å�եE��K,�g�Y����%"�OB���$"O�-S����<3.��7�IݱS�L��2j��X�S>�1M-��&K��\�-P�C�y�5�5>��m�b�g�$j�0�loFz!��k���kǐG��:��7�yo5�i4#�7?�pcH/M|�ć�/��TOOF�`=��z�kT�DP�y
5eJ曂���l�������O��u������ƿ������s��q_�L�Jl�y��*I��n�����\�������[MY���OJ�K.s 05�4�\����}*n���o���v�.܏���=a�d�K�����eZ��B�3�F������d,��q$)���A\	�9İ���pqn(����i���M7�9�O�H�"� �5�k�LhAM���9�b�U����2<8G4��T���C���ԫP@��ѥ�k�@��/_���K ���!d��Hd2����4�)�![%�w�����U����f�͹iR�w�;����eU�R\~֊��v��Uă�5S�o����dx�|(1.�.���RX��^� ȵ��`ܤ�V�a)��A��;�)Ĉ�VŊ����] ^��`���ɾ�	X�ǌ��}I�||8c�h�T�r�|�G���M�6s.iRMzm�"���"7m{����:�ޕ6CA����>�y�?���Gy鈕_�?���)?}�;F6m��6z��ˀq�̗��،�g��<�L8{�wS��b�=A�o���V�`ȩK���y�v4.-ۃ�
�'w��$�:R��^`�\t��Gus�>�.�˹�"2LSs�#$���LW���G*S�+��>�׻�6?���|k�'滆�}\h���������l���FEY����|ț��MHˤ�%��T�h�7��4�>�h�Z���6_��g��r1�8o�I�d}t�<YQ󿚳�P�$0p�`U���;!2���U�\
��Ip�x6V�S��B���d�'ż-/��%�Hl&>��d��v�-O���2���(�r��E/��	���o�P0I��Bc��4��x<ʐ��$�<\����P-���)"bB8���-R�m����%\�B�y�Z�K�NVG���	�����
���y�"��X�Q�0w���3��[ӌ� �7�Q�6,xq�=�VG߼~�3��4X22m?�[[ι g�I?*�����ƈK������+e���� Yk|s-[U���)��)�f�H������H�՛(ǆ�:$��K��_����Aim?���4��O127Y�	��gyv�X��5�!���Mg��Z���ɘ������Y^Ėq���%r��-3��S���@p��A�����sՔ��������P�(TC�.���vi���%a�c�ڭ����4�}������XFv
��wx�ZYY6\y=�i��FZ_�����z(��Z/����I�����f+�l�]+ s(�d��7c�S',� "�@đ���h�{�R��cۘ��?���L#�[��ltp2�J�rbXH2�;���(i13|!߆$��䊇�	��2���M��B��܋���Z��B!�^Wr����q�̱�8�4�΅UZ��&�j�h�&�1��NĊ�$���U�=�<U*���z
������Ur.{w�p?�2��`[ �M��z�E� �)�b���{�� �dp
���n����2f&�= p�ಘА��AG["�����<�\�>a>*v������6l$[�7P݄Kf6�0cU���0�Wz�#�������
����Y������@��z�)��V�P���U��`6CȄZ:F�e��֢b��C��ͮV�����_u�㈜�K|�sH��s%��%��j�+�A#��I|S�#�t@��%�
N(O��S��[[E�(XhG{A��^��H�؆�kD(0