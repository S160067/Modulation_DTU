��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����0� ����遼�6������"���#�{A���'j�Qj} �}xT	g��F����a��f��洜K%g==�Z���L1������bG����XB�k6T��w+F��3r1#�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>:��cG���Up�Y^����˚;���"J��+��sc��Y6�f$6�5&���z���������`dcR�+��b\�v���D���ղ:h�W��j����='�5Cq����7�r!��:l�6�Fo���_˪��k��LH�]!��0�H�c}��c��p��@]0��	$D��+�����7����ݯu�|��&��%'���潢(������,�Fh^��+��Z��[��b�i���j�=9�����M��Q������DRFw�G���J�s��2e9��X@4��b/�hp�� ��j�q\���&0%FF	x}�1�x�05F�̶\��6C�+gUA'�6�>���3�{EM��pfB��F�fv!��qb��@CÑ�Q�[��y��r�?#?8t\�m�Ǫ����������nV�|�|.����?q�a�S���P>8f;���$O��Qǈ:�V|}`G���lX/��ڛ�JV!�&P����[�I�

�X �?,'��@ݸq�F�&D�i�^� �	0l�{�L��hq�cB��	�	��K�-��SЩl�=�2���é(tKC��mA��jT�n>���!0��ٯw5�^L��r�yy-���@�Tk�ѽD��99[�I��j��&�S�7��NG8#��y�p#ҰӋ�m����*�g;ه	���0�t��b�g{�ɇ��R��:<�<�9_5���Ymѭ�Ʒn^Q�Q4A,D�L�ZJ��<8�@�15i�-�-�	Q�������X�Ǭ4Ԟ^\��K��g�_,���
H��:.�9E��Q;_�B�zT I�3�{o�� թ��΄:������@a���n��su���L�$�+�k��q\�@5bz��x�ǳ�e�h��@Q�t���8�tC��N��)�O�YH� �%N�'�M�yu�}�
(�����;�*��_ߎ���G0:%�3�}�~wui�i��#��7�]8��xZ�Ve��$�R�X�8.
+\���d�0!��R���#�.�2Es�� B�k�z��Q���[�&VO3��� �7,%���uw�.�㵬�Pz+��ׂgÑ7����*k+�"\g�[=5��cw.�62��L�x����w��1TZ��������<����+���yaf�7|Ǎ)9�"4�e� ��p�e��5���^��QI~��O_�?,�X��߀il���E��9��*1z��>	ǼzF��I���(��y���*0�n�ö2��#2fzDDu�BD�'�@����~R�&h Pm��}�6ZF�X�����6�P���̺E��dģ���:�ӹM����7��x�2�<Y�>/3�٣���ݡ�d�ǽ�l�w�Ǔ��I�^�8}�%&*~fZ�ɇ��D��cC�ڎ���w�vc۱ ���c ���32wk�ω+(R�L�^�L�
�=E%Ҳe���T;䊀�<��;�������p��Rxm���+���њ>�@�FO�'Gd����w��V����%�%�k������O�`��
��۝@\PXۈ����?&T��������x/4�#B)�T��2�P���	m[�"ب&t��j���`��O�N�5s��p�-���<��\	A�r,�)r���`ɶ%��ldCN��`�ڱ�~�-ZYex�Z�/t��<V~��Z#BQ�U�t@X2�[^�	0�^=
3�,�X�#�9��/��������=<��=�,j�/�5���/n���$�6�n��<�#�+L �k�L��j��͇i��d.l�j�X��&\1���8w-��0�dv���%	ok�s'zr���fs��s��U����6��g��J�g�|d �ٚ~~���d�>�(��Y"���F�;���Թ�<a'�;�bZ�N���ý��O�_�]�Fn��?	Yc���1{ ���w��,-��?%9�R�#B�5�«�(�}R��$�l���nr�X9==�Kܟ�mp�gl
���O>,#+�?˜f�0<�=zޓ�-B�89�`L�1x���q� �
�b�n���Z�q�|���k���%bD9�&-�8��z��JA:�_ ��n�^��ȁ�����*-��*��4��س��1heU_T�:�ĥ͋92��S ��S&zj�|Q�948S�l�� ���U�<>f�;AB��oIc��Zә1����^JKSn���ji��CV���;�JM�F�Ӿ��@�/�ކw,{#�h*g&"�;��-�̸��=�����JI:��_�EX-�j>͹��~~�����1�c�We%38C�oX���\�"]f��gL��'��}*d�������+�Q����I{S�6RN���5cn�L�n2�
�T@�@M���颍�~�sY�ɮ?�s ���J��(����!�X��Zm�F�4�H��B\����/�����Cs��k��T���݂%����sVb�KE�S)�9}"��ѩQ�HG�����|z��+���� �5��z]̜�o���r�^l�-�yȿL���S6�f����N�C����?�^rg.~Xɕ�b'<��?���s��
�!���i��%/(3T���ir�1���c0�uO�t�و��[A�����]�X
�I���گ��=?�?�4cB8��7,�s���[�+f�k�OO3�+݀Otx�����\��t?h�[y��q½n����?�B�蘚�V5��qq�4 ����2e�q���g�;]���b�[`�vZ��Z	����zM�2�f�<spR�����NV��:-Hc��1i�͝��;��W�&���	���E�FS �u�5��x�z�^"=G ����'~$~���x �R�X;T��tԩ��bÑܱ�2d����pL�ǅ��R���W{��7���"��7���B��5�Ho���⢚�`DU�)'�&4�z����k��}�.l�[r��k��G�'I�ե;Z��N��Q�Aڈ�#�[���m����*�Nw��ļ �du
�J45{����Y��N���A��3��_�ν��3E���&��p�qC[@�k�9�k~p�Vڱ�t��f�ju5�z
�nP�ܵK״����h�h\����� ���=-4�� R�ܱ6�H7A�<h%��W@P�,��?6OLy��\!�N��y���u�6�iE@xk$�c"^���;#���t:�6~޶�P�����ɽp��]����ҵP�)�H}��y�Wt�;�v���yG��3�?7�<��
wj��M<�$B�p1�]�AO�9��8�|�$p��V޷1�#�*��?{���)��Z �i:*f��*_B�v�k:��X��I���X��?�����}96�4���ޫٗK������&f��|:�G�Wc���9��z�H��yq�q���XW������U}'�������|��Ї�	%vCٻ�@�#��dC ��;�N�;�Sc˖�-]vgH��Y�N��ˑ�������!�����G>����zAq�� ��}e�j7�: �C����mͲ<?����)|k*^Y����l�0�FM j4������L��p���2Xj�$�kE�g3ܹ��t����s)$������d��?QmG�(*"��4��膚!;�t�h9��d]K��	 o{`�������>5Vm��ij��P?��,
pv�|��XSUn��'���U�Y���,�#)�Yt�%NVnYp�8��!}�"N\�;�d�Ȇ1s|���lL���'��bHic�#2d�;�׆�і~;o1: ��;Q=�W�0h��ɒ�S��k��akz��ꜟN\�Io_��Y�V���(�Z�3�ώ��C.��\�
J��������Y	+��R�31��cX6I���=�j
 �ZԬ��g�������A67F�e�P�Uc'��������O�.C����6��������W㮭F�����{i	�H
��9���f�;,�[�:�aL (�A��/sb��6}�rL���z�r���$�NWWa��0B����ч={0�}���b�������]iX*���c���Z�:O�qnS�V �l� �"��Gհܻ�����DA�=+
�\��E9y��8�����07�����}���B��@+cNm��_�գSt�eeM����CPF(�k^~�Z>�]h6@�����Z���<NC<Q/kA haT<ʾ���\w�Я����&6�<;g��]O5�ƹ�9m��6�	�U�,����Co�E��ه[�|EB%]7c��+A	����#�73㸥671�y�s���Lt/Ҝ�:o�+�zm�2��Ep`��0�hZ�\r@v�}��Y9
��ɱAj�s1�uB������\<�Z?:UW2�/����C��.U�X4��SN�(���^Wf���筶�6Nq�T �=j=sLY9���_��G�[1� C��l�WY�4�×��GA߽���/G��U�M�]�>o�aO��E�8�̤pM��W�[�%�C�3Ē����RA4�qf�ؽI�(Q�.L����⨩�(�C	�E�Z�@X�!�F�>CkG����h<U�B���RF����>�0��=�Ș��Oy�^����A��c�s颉��S+M6r��Q�.�ٔ1�DQ;�B�)�?�|�������j�mO8=;���L#�#�7��&
���T�S�LE;�y��-�c.�V%��] �r���NJ��,"��A����c?�OW-�޳5Mz�\�K��,�AY���Y�eMB�.NTXz��ȉ^�l�.y����;�Mjʺ�rE&8�[�ni+G�G�-��'	����Q��-�{�c#e�2�^�$	#j���*fi�v��2��#_�+�d&6����˟����LJP�}c���?�P�z��=w_V��k�k%i{�A$?�<������.+�R-�S��9�[(����k���צ�?��m���"���/ 1�u⹖ف���A4�۶_�����Taj}�0�5T�#��*��[�ܵ}����Ƙ�%Vн��Y$��B[6�t�k^��; D��fq�t�1�����xe��Y#=�ǃ��N `_%ҹ�zMۓ*��&�`�-��k��X$Cs� ʪ����Ʃ�;1A�	p*q~Mȹ���	�x7��րЄ9�^N�,�P�rj0E($���gB�⩌���ե=�t��_\���l�:gDR����A� J��dl�⛷{��DP��@9����~�$|ʧrt�����e[|&���u6X�[�ƻ�Ytw�:��r�.����ԮN�6�QP��Y�/�^*�X0�%����-�;ה�czV��@_�I`���4݉U��଒��~7�,h��Թ�wlY�H)X�\��l����nM�^��"s��]|�d�8�r��
q�QS��
����th�:L=-�.�u�����	�z�|ކ�ot�������4�]<�h>�dHL�4�O>W0$¸�Y7�.] 8�v(�|M:��ݖb���r���-�,���ͳ�Tc��bwKMx�Q��)8DJ6 u�lp�8�?ȫ8TB��V�kAKI��`�H%��Qe���H4�������%�y=הz y����=]\Ǯ`���

��F�}�=��M�i���Cr���#�M�\˴�aro*^����p�JL�������QzQKd��Ґ��I���5�t�Q%r����$��9��7�ݒg ��Mӂ�.��k��e��V;2^+v�����<P���p1츋/�a<��K�c��%�P�D�=T呅�)G�ݣ�ƌ^��>��>ُ� ���+�)�{�ɴy��ME�0m��Qa��C�����V*�]las	>�V�>_����Bٶ��˗ _b�PΈN�^�pm�����Q?��6IR�lu�+�d��Ѱy��^����_6yO�I�� ��Km�ដ�1��{�AD�_q���-��ϋ�A�y��z�*��y3;�&�vC<}�E��2E��N�p�B�sd�� n����&#��8��(�肯%��E�qH4k����uz�����⇀��A.��'������S�/�ej5�X�r~BˋoL�FyjoT����0��3&u���Y�xY>g�?�����LhVã������L���SPn@�>A�P��#�n�6�X�ᝤ7�,l�n�K$���� �/ޱJ�at�7W�)�g���]��q�"�:Bg��|f� v �x?pT�Ku�(�y�����Q�,{n$��(��6��9\/�C:�[����,K f9"�h-?����*�l�z�R�	�ȼ�'�MH];Ĝ���5�7����|ž��bt������W$	�}�*/��>殯�|2��H��v�E�a�$�/*7�P,>r�$�