��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���,���`�Q �����6�͍	),�6�md|_��n�x�"u������K �5owJh�E��qڑI9����%,%UEwf�x����;.�9��p3��,/�֤����"��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>c��mW���rJ(���/	���~J`2F�x���4W�0V�y��l]��X���8D�G$�ۻ��c��rk�E8o��W��z�����O�Q�F��?-_�䰹��Ny����o��:���l�,�:^�G���G��ta�`����k�
��^�0�4E,&��ݲ5)��اk<\�<�%����b$̛-�������M��!���p��Z����>D�~M\"��Փ�Kl?�j@wS����h�� �Aq����t�a�w}	qw���G�$M��t�n�^�lP)rO�%�'�CB�lpq'{E����6�,4s%��S�K���+��g���J���k)GVE�I�7��4�6��E#���'mಘ���3-=n2�ս[1���z̒-KO�H���-��rw�8�3�k2A@�8.)A�h�8k�P]b��(aG��^~��z&�%Qw��g� e�þ��Q4��/��8J�:���7��k�ڿ!Q�d���w�"��:�S�*� "a�~FG���<�y-+|���2�ǭ�l����n��}�e����3.y�U��M(<��4]��t�&�5U��f�ڲ�ثD������gZ�p�c��v��HGщ0�D���N�?*�B�U�����:���`�M�V�/��Yn�=��>P	���q����9tϻ�*�z>f�!V�]=`��6���¨�\�K�����@�i1\�`�����\W�Q�MXu���L Ud�%6�L�<�v���,��>]<�w�/5:��=L�D�( ��^��a�g��S[o���*?�)A����3�NhfH��?�;�ٛ"��'��:ÆMw��&t����H�ʓZ�s: �*I�9f#��U���qX{�%Ү?σ�C_G�H��$���@���+A��pX�� �z���顇�I�Æ]>�n������I�	=r��W�î�m��0�mju�9�q3���N�V�7<�x��h��A2�����ot9����{��`7�vnm�Ȯ���S���تUF����
�Ě��PR[R���0�^�����tH��v��y�Q'�SxƟ_	�<�#�FA*U��UJ�1'i=a����LEb �"Om�]��{	���.�C��j

Z`�:�\���P��!� �bp�~�BGHׅ���1�R�11G�h�jmM�m�0z�]9�n��4[ydcw*T�!ըX:!;��tހ��P/�٤��(�@P�����{�g�9_մ���x���]�A<��F��J�*<!�VR��֠ܐ�T���]H0��|SΊ�䫎���,i��������C�����;�N��	^o��n�_�t��h>'5A�I	�nAd0��O�cv�VFv r�R��H,oN�{��1ƪ���訃>JKt^�n��9��Qg\��i7*B��(*Q�q�Rw��:fSF[|d&9��[?�'��'E����9>���ݒᶷI�<��c����QV���xuŃ�`�={�$8����H��F��qL�����"�z���8O�B7LSg)��~@�
V�wa�~a.| �}������]����;�B��M-k�4ԴJ�:�+ýѬ�[�Kaa��{&^ݮ1)���$�v�؎��� #��&��w�,c�I��&fm��5�O.�����P�14�É;���+�C�W��;�E\�xZ�!(vm0�]���� ��� �F�B#a^JOehDf��dC9������^鎾����)������0#���%�f�Ia�y��;�?��3�����8�+)����r/�²�SUlЂ^d��<�S?\�V�?_&;�QL�/4�P8�\"'�++�/+M|�F�V��	��Y�X=7@��`Q����x8��+Q���!1q��X�u�%(��xi��.�l�٘���kI�	�,f��
�rK�S��p ]��`�
V��%X|:���6��A�iY�@�	�3��0�y�4�ձ`�rG�ԗo��EH�x�)�^�y�J�y�]�(�$�]і(3�Gk���0��\F/<��j3�y-�Ë�����}�lO�7���0x5�Cv'ޏ_"����]6I���y7!����k����M+AX����Ra�k�����S�����a�JC���a�ƻ�����+���ss�27̅?E���'����@��H\.����=])7�����yV%	'嗽:��u���c�Ƴ��V��rI&��n�f�K�KS��[��Y�ՎO�9T�=��Cx��/�wl������u7�Ѡ"�X���-��GT?��SO˜���Pn<̜�|YI�F����rdlc��m��y�f�ي=����~���
��X^a�q���cA�~��٬���@i����6�o�T������5�S,T�띛��U�����z��f���T�Ȅ͖&�*�R�v' ���F�`7�B<�-��e���`DC�}�8�Eɷ���́�_%�$d���l�$�p=ݑQ������μ'}%t�ڌ�c]��貇��M�n�����?��k@�n)�c�i�\MA:T�䳡���riQc����{|e�C�����5�0{D����\�(�^%X�y��|ˡzd$�(��"B�cu���,���-��c�����L]ɩ���l�#�:���Ь)үr�Ӓ�!�Ε���,��VEZ���j�!Gٜ�~M��ӣr��g���-�L��Q�s���?f�)�����"1{�51��=)Y�R"�l���_��O+�ޮT;��`�<3�@�7�#>�.(���9k �����S�$�k��
}x�;�5�KLRE�v)��>q@��`׉lVbm��,8cY	m��-[��Db���J��S}�*�̯n�v|w��O��5 '�tuC�CoM�k����$C�<y&A�º/N��E���t��̣ޞ�j�t��2����U_� ��Ŵ��Q�ً�	V��']ձ4N%�f~�_�����,O�ȸUH;.V�[?��<I�j:���.F2��Vs�O�� %�zhl|�_.H~�=���d`��Q����r��+Fg�(gk�l��a�<��p�?M t��W(d�������Jv�3A����8��+Ḙ?�b��AӹC���4��i�T�����͍כ.3���ܦAn����Xҭ��D��i�S�6�};H�6H���<"�o�,P�+l��~]���s1�'��me�W�ۤ@�1g�	UD�����
��U�*]_L��	hy-G����t-\[�	�Ku
���3��	�$>k�\�;A�`���dZ���&X��O.*�f"B�Ij2'��Y��%ȴ�p+��0ۆ���Tp1����Է�!��R=������$�uv5�ݡ7��q4X+d��