��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����0� ����遼�6������"���#�{A���'j�Qj} �}xT	g��F����a��f��洜K%g==�Z���L1������bG����XB�k6T��w+F��3r1#�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ�A�O�c9b��2���j�:��HA��?�\/��q�k��#W_�0����J杦�&���£mj��̟鬶�Pf�s5��q�Җh.�k�/��HJGS!]$�y�}�t+��`lJ�g����?u����pXp��8PR	�Z�,&�gtL�@L�Rbӑ�������Dxb�2�Tt�����{'j�~:9$>�]��H�� L�|���SV;��o��z�.y��o��s̅�0��y�h��j�4?�l�n�����h��^�V�F��b_5uV���r~>�;�`W��@Q�z����6?C�Vܒp;�4Y�A��4퐣 ���i���h���J,���d�(��`�i[�	�X*�a�d#��/�`r	�ء-\Lv��ɾ
K0��r�:U�i:��S���wh�vP D����u��zB���Q}�#��`7}d$E'$h+�LD!���j{K��ϖ�"8Acf�%A��3؂q��L���pjsմ1/��W�Uqp�ʲ� 0�j?������=�H�+�W0��`�� �h�.LN2��=ԕ7����ݬ=d���L5�X�»��I9�&�U�����Ɇ��AQqr�VJ�>�9Y3'��(��*K�a�
C�uj4�����&1g�3�jVd��m������Q���X�و�b�	���_�3��07Ӷ�NO���y7�;�����
pa��{q))���ލ����T�����lI���4'^��U	�\&w���E�� _�xF/�|��[jMVb�����liZ/v#ki��- |-_sw�2� �4�)�w,rY�^���&��̧^�l�p�]�6`�ҥx�u�]ɃH繎X�YO]�5����-�5����$p��ƌ%�Ս�����'H;�WF3�`�uS��nx1vK����h�薬��:�2�������T�k��U,��������kcƭy�]�zݪr�e���0�d~(�A�A��-2EB�.����rJ|�����t4]Q,,�G�th��2��B�^P|*Hժ���)Mb������X��aX'�׳���F��j��o����/��C���G�9esx�o��Wߠb<� 3N�p��P����~��m�,hGrHX��+}�Ws��a:���,�0���.�9D���;JoԵ�4,�ӝ/�u�5�Q��WR�9ݽnA<���[����1\���e��ui��&��}�ɶwwVW=�o�y
M�M|n�;u喔l$|�/�g�FWzO�l	��`W�\'��h|�}��P�tԂ�n"\�m��$m�x�����BA��d�]C�{Nq�τ>W�+z��bb�t����j�$QT1ř���g�V��l��)��[5	�y��A*U�p�ڙ%'��0BP�֧��"��-��~�E�2�A.w����`����c���$cdhz0�4f9� ��Q��:	pR[Li�v�j��vv/|t{<!�Ȃ��xZ�`����^Չ�Gi�61�4��8��XQ�V��0��h`��V����#�J��m�� �Z���PiS��е�i_)�9��l�������I"�T Z'C��t:`c%T�H�(�"aƀ�K?o	Mp)k�G��4Ck{����ce��4v<7�]�j���8։@��F�[%�NAr�>h���K���-�NHO��J
Y±��hF|�
^�,�{;�a�ŅZ�G>H59�":�tu�]<pf��0"�	t[{v�j# w��6G�^�W�j���8��$ھϾ	��ش*y�`}Ԉ,���+��k@�>��������Y�w�Ƭ�-*�b��YО����ۡڳ,�?�k]���ޕ��#o����n
��ٸ39�CSt�E˨�AQ�ALJ�{VFm����9��Z��80G9v��V�La�<���LoW6�v��xH���,��\oU��H]c�w�z��ц��}�ݑ��Г�_�|~f�ܚ����:Cn#�Nk���D��K-�'����A��=��9��e�ET�HC,��� ��f��#��
	�T�a�4hGoą�M斚�]�m5��}���{).������R	(X��AڛB��܊��=҆r%}���N=p	��`�z�m��g{�쥈�����a�Ĥ�X\I4��H)�,���'�Ck'�Of�1� �� Q���@���.oF���Oxel���O�#h x���W�&�o@/�� N��2�����{(���A��ĮqB�]iD��a�G�=��^=��������6�6���P����qЈ�4�H���6
�����8�.i0N�H
tı��zl����7r�ῂh������Gm���F�&I	��o�l��S���4�N*�FQ�G��=9�A��R	���!��!t�{k�&&h�u�ch�XWH��W�V�qA|��O�g�����@,�'~�=`��è�(L���=Ğ�]�(�U��d8�s:UA�K.�C~��e��^�<����� ?|�e�mBo��_��v��א�4�[��� '`D�-����Q���WB�����@!4/��̭܊������_�'+�U�)�g�]�<zC���ݮO��n�/�1<�C��3�zL�{ T������F`�(��I1��@�_�ncB@Yi5οƂ��s����b���<�j�2�i�|������A�@�V�FN�ZN��X;����Cʇ���7�`�f�Dak�m�9�U��r�����<��|U���ѹ�����Ma�ɨ'P} �a����)Q,�X�ė��h�ܜ�*���Q��=�����~k�*l9�?ڕ$���}�*�:=y�@�vϓ_���Z.��[����/�3(*#⺻�P�;T풺S��1��7T��P����0�lU=E��	<�B}�)��5�z)\���*�{�+(m�B���:�up�e7��D��K4��.�0�P�?O8��\b����������+̏�-���X��� ��W���k��ni�w���~����x��L�ZO��*����Q����ӻ�r�#�N?">y��vJR�Cu�e�S�{w���cw bQ���m1�ZD�&Hȩ�H���0)r�|�,�?�KJ��Eq������&Dd$l7��^N+o��t��:�:��Y��d��\)3r���O#`��B�����ވ=7Iĺl�C��s5�$��c�	a����ϼ[��ްA�,	�
T% -���Z#_�GJkZ��C�����u�����l��կ�L%�O�N�'n%�VxX�^���Q,@V|sڟ;�R�	.����������u���.h�nA��v�̐����64 �5��!l�}e5�ƇZ��VB��L9>gy��]Yd������Rw�$��T槃�Ph��6�B=�S7O*:�6��\�^�U���Q.�I�o��l�̣i*�h�{���#%�Cy
_�V>�M�������zs?л{��W��`�^��<��)��J���N:S�*v�$�.�b3^FU`"�A�CB�U���j�Q�����)-(� WBE[>���9�_�v�E"��f��\g�B5u�>�[�<[�c#��a���I>[��8@nm�Y�+z���9�i����%|^1W�@-|݁!�@����T#�3T�<����$�j�@:ɳ�u��eF��='؄Ҏa���u�s��A+����V��g�_m M���_Vba~@n�U�f�U�CL{t��4�����jY	A-�\-$Py���*�L4#�2���G�&���A3da�{?+f?���y��N�q�*���PU~�N&Q��� �D"��z^�_�k�����fC��_=�ʎ]��ӊ8*�_�� ���-������9~��,		��Z��}l!�XT�Щ�(�Iu���O�:rN��j7-�-�a��q|4�־�����=��˹��]��-_א��ݲ-��Z�ŝ#e�����+�SsR��Fsg]L��aq@2F��C�K��WZ�2g7��Yf~H�Dǡ��M�W;�s9k�V@��z�=�g��c�'��gr���D�a�N��+�>0,��.k@Ԓ>�Y�X��l�$�Ӕz/5��/�V�R������'=w�v�STN)T����=�����\Z��	Jݫy��Q�����0�k��|;7'[0�{�S�.���t��!8���M*���>�cHW���g�N�����BqiR�n���aP�#�VX�'E�ʎ̏��0_����"�%�/��BP8ɣv��\�(#l��5��k*\h�a[�?j%I���(�8��isL���d���3%M{���fkNB��� �[FA�.dy����R߳/N�0��*�\���$�k��N�h]I���we���YN�b�9�Ғ�?Q�y���帹h� �4 �|��z�4H�QX��v�<�ǎ�e�w�pP�"p
$7O�T�ފ��Fl��w��ʳl��ټ 2����Os�~���JY1Til��3>�(�w�����[�9L���e:Uo[�D�qҡR�<,�&w��#�)l���D�a���śn���jlp7AC�W��P)
��;ؕ��w�����s��+����Ϳ�GB�d���*�3M��Xm�>����?T��U� y�^�ɋ)J�)K��+���/��	S�L�u5oꠁ9��+�c)3��q�[����uȖKJG��x{j�����HF4�gF�fn��(P��4���5("�=�bXص���r�2[�G��i[�����kj���۵*��o�&�%*��o�1B�����X�;H��N�����M:��@ʭ�Ms.tc)����H�t{�?~�\ҤK%1�X�X I m��AY��k�[��ŗ���?���k
;=��r7�k��k�OF���x(�E�f[�󲢂�m�4� �D c�D�+�wGy��;� P~YH"��:�����(-�ٺR���Q�j�!A�x����o�_��q&�G���mE��A��Y��P�����&O��d������)�B1b�>i�{�)����?.�X����ϗ���,rP8�����]��o2ߊ|h�ٴ�wV�M��@���a����/Z���*nbyZ�����C돍�5����������>�"��R��2o���r.e�	H�~�?���N\w�;Q�������8�R+�ձ�aܗf�H�������u�	�LX�ޑ��c2���l���%/�-%[p�8�=#�bn_�A�O^G��~��K��B"&(�݇�$.�u�}��	�Y�����n��x�ۼ2۸��vˠ��-Gg���3�j<e��b�肕���_�}
?�dS��qZ#(n��˾�S��q:c5-OD��'����ܦ7�-�;�,�|�����ʱ'2���+�Ψx�#�_�4M�9u
C_�f�h�.^N�NČJ$RsK�n���4��U��ZA�8|
Nt9C�K��8�e#�\��B��`�b7/�d�&���_�&
J� Xr�����{�B �@�x%��b����X8v�L��`�C����m�S_�KT�g�]��,j�}*g �"�3跉`�c�	C�@��XUp�u����l�bn���N.��@�W��Oe��c!P�%�Rx�LnЇ�x������;�ӵ�w�p���7F��o�_�Y#�� )/�������h��M���/m2�"I[	��;�}�,�B����"�N����"FУ�lQ�'�����C��<�g��1�6�M�JO��K�]>|S�8�o@QW2��|�h��\���hh�����Z���2��?Ò.eg�n��]N�J��'t��2�78�vG���;�'2���s��D4z������(i����Qq����G��A(@z3d_�c��~�����sl"�ߗ/�R�o�}��2Ж��d�����L������t(�����ɨ�os�1eM�OF��WJ	�	/l�Dԡc��o>�{$����6)�
j�e$��Occ�x�3�3zDʅ���;`�v�lz��NrE �Q;��o���|��(���I����0�g���M��A�1W/b�w�*LW�&�]'v���8Nْ���5b��c���x:�`�
.<�%�PjR���(�yHX�����΍'|R���� 8-2@�^lN@�*���a;s�����ͩfU��ǖX��kX�S�%s�\��)�n�j�P}���-W�k�1qO>��>ؓ�R��c����r:��eV5�M��O{�����dE#�ٛ���	[�f����<s�,�/eN���4�I&خY�e-��f,i���.x<�ښ��C��#Ђ?�]ri]�����AC@4=c(���V昺A<�e������Y��I��DU�ɘ,O����y	���â���T�[����JC���1�&�g���')�|en�9w�HX���[8Έ��}Sv=/%�g���߂$�J�9�g�O1�F=�n����nh4e��u�!��
�0E�oX:����>�9Ǜ��w��e�i�(�[jȾ�J���Gm�5��
uv�� J�)�Jx�T��;��$sY����g$Lhr�'9��D|���ͩHW-!�n\�o(P��|40���ZT�O���6��؊���8�}����KEi��ک��]UA�����n�I6�6Փ'A[H�V�|4��{�4���f��Ƹ����A�Q��:"���IE5�u�`%p���-$�0�3��'L��=z�]d��X�G�F����f^]U�� ���9�4�c�a^��p��$���-��Q�g,���ͅZ�I��ѯ�G����,�C�u�|Q�dD?M���v�EP��t�ҕ���aﵑ�`B���Q�d"�E�;�]�)�3Y�(W�SW�ϾV��~�3>	�3�����R�)u~�,��ک��d����'�|q���"O�Z����Gi�\���=��F�4[�Kg^J4o�$�0/~w����i*K>��x� �φƬ#6=�\�|)���b\�(}=eG�����]z�r'���]�fc�Nh:"���{mq=w�i��V���q��L���p���׍��?��¤���7TE���f.)�ؼup��6�z����*��#�ơ�?�Њ]�MXN/��!�?ۢ�V�6���1�/y�Ś�R>x z���R����'F��s�RX,Z]qI�&��gp��ˡ�	�T�}�{Q<�8���\dh
-�d����3䦦3L��ZP��#�5���/�rX��(N�V1吪���jä�Є�mn;Xs�G��r�@W������t}�3��}�����l?�0��C��O�"�(�͊@r6�+�
�))���}�TfN�7��Q�h���=��?��hv_B>v����On�����E�I�^,�xƬ����l�l�]!
��dp��-�I��_�Ĕ�c�$�P9�����tx]��������ٙ)�A�8�|��@���<��J���}0�XU��t�}UOʜ�%�w��؃��,�Gm��6ȞW_z?Ry	?r�F�J_q���ǉځ��i�`�&뙫�c��ra�=�q�_�ҫ*��F^��%���7��;�-�4���t�g�_�7���,K�Ǫ���LB��C��@$���h���CA��(?���U�;���_ך]��t��2�V���X�,�a�1U��L_!�S���`�(�Gy��9������b:f>��v�m�DB�	ޙv���P�ċ3U��:�S�VZ�g��3Q<�W��n�5`WMc�`	�t�H�g
����P�F[��/�C)A�S��}z{V�N8-m���.������'v��o�f�����7����aE��@�x�����n!v�1�-$:}��p����
Qa,��&I�	��mkg��?hH(���U�>�,(�:̾N�<�]��fQɻ'K����ܱ:�f��3��#�߭w�_y�>H�b�&�����D�'6)�a9������WD���L�}���������:��A����hgce�w�y6+�Nn�>B���&`*���L~h�=����~Řy���k�$�	JS����A3�/K�4Nvn�����l�9n #o�8�|�k�h�����{z��n?b���	Z�*�X�:ø�u__B(ǁS��4T��V��M{�_�Tu��v۠Ͷ ���|�	�:�q��8�p�e&O�����f��[>�q���l��G:Z���Q�M:j�Ãmѽ�{�OD��щ�Y�嗏�� ��@����$�:i�"`�㍠պ����j�3�1�n�>������a������w��%��^:)��TcAH'S���a����ٲ���S��d7���Mó!�sթ���e����`�:��U�|eN_w�w�\�B�r@5&�з�� �����{������3{EOwSO�(��4��3օ� )&9?�����Qc��)E�9�#��#��d�.:�G������:}��d��M����m��Ǫ�o��V�2Ŧ_�e1�'����"7a�C��@��.�x�51��Npyr���w��:�`��S��w�;ĕ��� )D� � �o���JԸ��w��P������TT��K���!���*|���>"�8S�Z�g�B�_=3���G�~N(3�ʭy.o��~�����q��ٖ��1�>�^]6^]*�`�wu쫻��ƾ��I�Cfأ罺�EDl�{��u/�r"�.W}�MA7��ߚ�[I
�I��Ν�ͳ�.D�}'Gl�aȄ"r��Fnw��-˃vU�n��P���aUu�*y%��tK%�<q���.��T~�g�n��^�tK���EAec`ʺ�L�v���ȺWi�9�G�g6뵆4z�;��,T�fJ���p�������Qr����qVw�*�F�/�	�u��eƂ�,����z�ѱH��
�ķ٬ ���bU�3B0��Dq�)�, u��	f�M�e-R�)����>�U4�M*c#�e.&�E[e&t��+����pl�6驅~��D��ȇp�/��]�Bn�?�/������Q2r�g��G����zM�l �;��񵦻jh����E���܃C�<Yx�0����~��e��L�7;p�~�m�·��kmb����a�8F�J�Q��'&���%;o��T��~IF�L�zz�!K�Ec��SWO���7���4m�Vy��#�^�G�)�������_\��--��1��ޮ����r�l:c�O��k�Y���:2��X�����`".zEP����x(���7"':W-д�<�"M�}�$F|��t��w^~����+nh⇨L����a6,$�M�����z/���j���r��	���������t�)��^�9���
ӼU3I�>�N��f�'UPTy�a4_:�O�n)b�!�Ԙd��M����P�NE_�w��/�yM�0�נ4&#�u�,�v�m���i���ꐽ�<�O>2Z�y(��01!�K.�l��3�|f}`����xݳ��\P�dS�s�e��b(�ŋ����7u=�����7M��:6���e��kF�ۺ�U��	�I�װ/�Q�������`�����;�l&Y-?���?m_|6�y ]*#�AH5�bf�d~49���m�T�=�X $��@� W4��:�����R������T
J3#�L�=�^�}�g��P,��!�|\�#.]�]����G�����߬TLԛ<kY�3{s�#����;8��jo l�����A��Ob��9B��AJ~�򋊟\�˯��
���.�\�+,M��v��~�^�&���6��Ha�큠?�X�sҳ�*�%ʳ"�e
a�ܘ��2�<��xZD��Ĩ���\�m뛞P�����-$Di#�n��>H���������������u1SD-���B�����٤�?S���!c��v�1�����͛bi�'��[��e昜�>��eL���q^�����Ol���- �� � YGf�|��2�H�7Ruк���J���Ñ��[�b|jC.vC��C�74�����J�9�zn�B$F�l��5 �q���I���l�ڧ�맮@�ڤc�R�@^E�]X6�����k�;^�:�����9b�۲o��/P��{����K��9�D� �E����G,D��ՙ�v\��]<�e#��Q�c�U91�����h!l��Cb5���UT���R�ލڀ$���`�����j
��mcد�?j����k��~�������Մ�-RZ��J?^�{����Y7� ��dslNu	���{�9ꐔ���è(&��(f��Ԍ��pd��<urvZ,��5���
68�`�d0�.s;��*F@���nF��_�bQ91x���$Puϳ�m���:��d@�:|�	��4%r����(�-�>�D!:����Y�l�ǵ��Z&�~h��$�H�鄌���Zr�ɘo�(�ȑr�$�F�0l6�?�a��3��2B��n��($�	р[SrJ���>s~��N2@��j�'�U����L��\�f[�Z��8�8���;wEF������X���E�g�B�FGY$�{�kܸ�+2g�� ��ǥR�&n62I���m��%#�-��I�yR�Oĳ��
��3�z����׎�z	�l�w5"Q��Z���9]�W�O��'���� aE��𥐍������I��)�?����⍉'�Ѝ����ڤ��ZfE������� !�J���F�%DN� �����Tل��ے��Ջ��!�f�6�h���-��@4p%`�X����bfǑ�**�E���)?>�}ĝ'��촵=��{���_�H}�3��� �*�^���+���
@UB���2U%˺d���	U�S��3|��|�H�o�ǚ.��9qح��ĽJS��Q�Mh<XWW"z��[�3"-����>�$�t�-��Z�-ͫl�Ցm2�{�)���CA��N���/8�m�O�\T��Ru����	Z�\e<
�Ղ��LXK�t���R��xd�t@:���t�[&a&"VU�d��+ߧ���-���j��? ��ա^�cs'5nF��wȃ��o�6��c+$B��?}��_�C<H�+Ȇ����w��w޸��I4�~��"=y��e�x,D�	�$i:���+��ؽ�	�m���,L�t{�%K��߀�J~S� �0�(�Cp�1_H�C��	�'��