��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����0� ����遼�6������"���#�{A���'j�Qj} �}xT	g��F����a��f��洜K%g==�Z���L1������bG����XB�k6T��w+F��3r1#�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htdʮz_�0�`��@�[D˂8��k�ľF�n�Ԥ��r�τ�u�&&����\l&�$������<H�����}�ƌRS>�(B-~�� ��ڣ�9#M��c��&��C:��p�@n��7Eͩ�4�.)DQ�\w�:d豲:���b!<M8���ZZ't���s�q���(Ӆ�>����s>����P���Jr����Nb�Ao�\���D>N�1lH����+������^45��(l!�,X^����vqeW	iI�M�ж��v�����犰��}w�>V���jǨ�mG����="�fU�瘘@�,����� fH��KUb���ϥv�����2�#�9ɠ��qk�.*̫�׏��͊(�<2�at'u�"朎�����w�
l)���Ѽ�!]�˞YK�H�[u!�3��X�U�4�1z�R���@�v'<yv3Xٜ�wm���ȧ�Y7��m�<��.������c3�v-�ek='����R,�զp�rw�BM&&�;6��c�����f�����%�\e.ac^GS)v�e|�Ѡ�⭷���<��x4:�ʧ�?5�!��U���;e4Cw�>�,S�X����/6?ƛ���&}	JCZE�����t�G����Ěg�ә�Ep��ݹ���e�(����C�]u���]�~�8N�DT����R�.��S�w0�E����g�;��{A���bݩ�oeZw{mk8�O�uw'�X�7Z�Ο�C�D�*�Yoñ�R�2,h���(�==��=�� ��5�7i?������dY��ɝ
�,8^�6ґ�B&�ZG.A��;4Y�,�M��~�e��>�( �kX�B�����aϞ��B)M����qo0���5S������
d��GgI�;i��jy�znG�lS��,��3�E�A����;�s6Di�CuI,m��߼F�����K��3�H�C��~)�9\RL�&}C<��ڐ�"�oI`޿\c�ALQKJ��x�XOlj�������oQ�N�Y��>�D�ࡋOR�@|�]������:Ж��d�ں�LY�r�6�2�)��u�sH�/8��A�����������EB{����o�o�	ʌBpt[��:J�,���(��o/I]]��[6$rsG��F�fZ^I�c��-�-|��?�$�K�<cm���a%��M�M>U��r?[&b�H�2ųI�!Ë�WX��Ibڼo	h3ߒ��˃�1�!~`�3�o�1���D�?*^uܩ��s< F��s6�*��l�Q!R�Wņ����:�~�}��Y�i���U��"�,S��ܾ����0���n2���I]z��8��D���t�"��̓ �4�)l��h
�X���VMN���d�5L/ky{æ�XVm�u�J$��LFGP�B�rd%��7�>�)-���o���j��ʞĽ
-z���� \Q�5,��n�tA�ì��R�&��b�C#Fv�L`ˍWY��i�+�*�;faC����H>����c.a ���<����t��6O���x�>R�/��O�ť�ȗ0i�+fw�}�+��X~i-���
�pL�����sG
;X�����q�x�����ΈQz
��e�p�`��s�v�D�m�'����x��8��d�ԘK�W���� `/��'p��-�'9��B��'�w�)d���-�T-���టhm��h�b�Z�TgZ}����˽����O>�'��>5pC�kβՏ�O��������s?����E�X.U:�J�=?�坣s���W�ZL,����g�k��g�y	�đ���������<����~�%�$%�f��[���� 
JG~!��l��-���n�ARzHκ˾�<=^��1]q�U�>q ����G�o%����i�ϯ-��^c�Vw���XQ]������o
eb�oR���M2�6�_kZ,,�k�a�;���#�izI�P���AT-�W� ����t�kk�$��*ƟQ$�_| V�c�T�O�$���*��?!�S>wJ�7��U��(���4���	��<�w#s���M��:��w9&����[b�#`��� l����;w;���.�]�>�oPz)\)�Ur�=4B��h:��y���O zl�����'vL�n&gS��%��	�u�dͪ�+N�T�F�=��jN\l�"��@��b_�Hy������}��b}�a;
>@�G�n�5��:Y�K��f�@��9q��&�ĞJ����	�G�k�qg2��8��_wX�.��VO�)%uu�M����-��'������͐Q��V����z�r������c�Ѩ��_�#��U�(���&�:�EhY�0�?��,	�	o�����$[tnPn1O�ÍW�]�W��ȉ�����A��!�����*�T��Ϳ�|ũO;���Q$�����3U���c��E�k��k�]j�����o���"q"I�t���=f�^��z�VU��ǘgPp�� �+;�̑�;����$�Ay\�@��Tj�U����k0��ǧ�jy}t���:S��3gwRO�񺓒��ПL�M��ߘ����c�	��D�(J4l��A�n�y;�{���U%���}+�a�<��W1L���J�%�υ�P��O Kwdc���R�R~� ���/����m��Q0�2D��m�8~���J2�a���rLВ��Y�C��q��B��3]:���ʌ
�<(L-����v�+K��i����%%?�ޫι��V����:􃹪(���w�C]��E�Ӏ 
�%K��"6@`���D��	V� �b!��x�����փ��QG'�K�b������\Ʃ�Jp�@���L����YfДL�@�%2�?�,Ӥ\�;$:�>���vH���L U/R6����<Hβu�b�<�i�
��ȵc0��\u�����_��yǖ&)){qA�����đF�Q�a��1��V[�A�U�����&�&�zBӪ:��pM�}e�\�*2�	���h%WZ4�P�%6w�t�5���5[�O�&�p�AWG�x�ʮ��t@I�%X��� gz��Y{V6��2�U�,���%	
J��֐0A�>�#t�f|��Ε��z=~��*�<ߦ��H7lR�gs���ۆT���V�<_N0x|T��T���:�A�w�D�G),>@ %Ю����P���XD��˲�)i�).�-�(y�r�sۏU���y�n�0g�@nk� ́�G�1?a��2� ��n4T��\8���e��f|BU��L�\e^�ʖ�$W