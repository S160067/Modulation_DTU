��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����0� ����遼�6������"���#�{A���'j�Qj} �}xT	g��F����a��f��洜K%g==�Z���L1������bG����XB�k6T��w+F��3r1#�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�O�p7��V�ӵ�c�g�g��)n�4��'8������$�qg|����3e-Ȳ�w�BQ�Q�w��.��A_�� �����7�j.k*
�? 
��#������0O֭J9RQ����wY��"�Cm&�Wr�+æ�/���4�ȜP%����dō;-q�������0��j��uў�������<���KD{�-��ϓ��V�wYB��,Uc�+6��n�~j��\��8/�hS-��)<3�CG��Dumy���mb��8:)(���T%�SO�4�39=MYx3WG/��ǐ����IGP(�~���f���K�_s��n�������;��޸47�J����K��a�L5�|�:e����4#��B��@ڱ7p����!��!1�J	�qV�N���K��i��0H  R{Z#捦%��l�d���R0@��A�f㶃��l�;���Sj�(�a�AyMm���2	9:�����*l�D�g/6C��@�l,2L<߽�V��
�`���W�I2H���I�v��P�]�a�Vu �ݙۥˤ���h"��L�<)K�a7�O�~�����N�v{B�z�{h��a��⣇3� 9�ą7�o/���`_\�����+�c�}���ϻ��Mq�0��2�!ҽT����h{��7f���[0:EhyQ�Y���s%>�4?9��!N��E>��y��5R�*���5�ed'��h�K6���Іz��.�FM�a
�0�L�S�����m5fX_%���_��Ʌ�]��3��{�	�e��Ҝ�6���g���� f�J���
̐��`�k��yjg�/��
���j��x���&wf6 Td�|�ce�Nj�D�Mi�(������ƭ��ٜ�qGU�I��tN�t�ؗ�;���pp~���?f�&�M�C�pu8�܌ ly-$M�6MĻ����9�\b�/Ƀ�6ن#��C�@'��y�i�F�`aB>������A�`���d�]GX�A�rs���^����a�ʔqۆ���5/p{1q͉&=�D�~V©���rn��A��#:@��!��c���E@)n��2B�0y���;������Ͷ1*���Ax��[�mHH����-XX�	h�5"�-4�?���w�2�P��na�uF�m��YTopհ��"u�p��P?�=@�(4��X�.��+��!K]_��.��g��#�)���dͳ�
��63l�׮��o�x�T�M�\�4V��R%�zX��YB8�gL��8|n�([�)
\rb`����,I2����~�m*p��>�|�D�KR����\9
�D��E���bX���v��Q��$��@���6�eB�m�w2.���mՒ`��|(�9��Z��8e�gɪ�2����Y���T��Pc'����D�9"(� ������90��.j�� 	Ky�h�=����:�4+��`;�,�b��QZο ��6���ܵ4N�H�����TD'��V�z*���,���xe ���ڳ�U���)R$��+J�n�� {Q䰛� :�I�$\ d�J_�v,sm&n@�.����ha\*e���^��2@+R/.�s/1�R�t_e@`8zի�d��r0��g�<�$�Z��-����E��[�f瀄�2��D��^�T9T�n�9���K����6g�tf�(���G�+�����k_��:�˚S`�n�����7Ă�\s�Z��� �J��V�`M4�����.��):�X���u+2��@	�b/�3�VYTG��<�й3d���mp��^h�C�aW���|s����H.L �I^��=m���2�5
�*�+��cXB���gc*(K����q���8�y:��; h�+���4�#�
z�(�`�]I>���=�i-�J�$�@b/��e���G"ϸгB�jA�nٳا�v� ��z��{Lf%G;S<����F,8b�Ҷ�Ԭ�n>+�5x/�^�Z�D��!�j̖��u�Pa���+����F���)�.�iG��v�L:����Scq�43�3�������d��y(ܫ����o!m��9�s��;(�L�|pM6X�Z��S���B4���Nߑ1:d�O������`Ýe��7;���q�[�̿<|��,g1	��ɨn'�,�����2��k�N�`�q��`}���*����h�MV�$1�ص�W*�~1Az����s�%Jm�SjX�T%��8��}S��X��w���g��OE�w��yz��:O�D��A"����o ]_� �W���6���߀�I�	��>@�kjsE��s�������C&�˼���4K��EL��a��
 �qf���d���&��Π�L��nJ��d�h+C�^T�8m=�y����xOT�93�i�D�>��^�/7D��p��8��;C�[���G^I/*��ⓑPX�^�O�����K��T���������������s1��	ٛBo�f������R;��C�Ȕ������=sr̖���V�D��m��(�>�jfL܍qL#�=k��-��0��������b���ƨ?�=$T�>b��J�{Y�R�V�N4�����'9�O��~�O�{�*�aD��Y���5�A8�ѧ�j�K��� r0�ҩ��7b�M"�,Ôf(`��nR��Bʖ"�����$���I��{�2}\��R4|���77�����>�c>���P�vA�|�s����1���@#��8�WS(�{�RYZ������-Q=����Q	JV�Hd
m
�~m?�h�+��Lx`<�K)�?����E0��e��(�U�9���p�A^$4c��z%y�A!\���I2qP�-jY���^f���?�3t��{���ʝ�n�!5/���P�<%����g���YͳW�+�eyol�=T/Zt}�:S=�?�'�Ȭ�j���jxr�W�i�'��C��EI�l���ł�
�7rY���)�&+'�V0���al�?&�p�Lp�d�����?���o�p�z�i����J��O���d��GzϏZ-��B�ۣ�,�����ݾ��'x�Oq���ɸ�3VV0��m�:��q�Q���p<>�fɨ�$�����Vt1o2�ŀ	�<���O@�2dg��ް�e~Z/��Tڊ����[���{��D�B7����it�Bj��à�@ІN��6`3eHÁ���;�	���!NU��6-�k�J
�0Y���{�;���U^{=�ܒ`�DZ��F?�I��M�t��V��J����BT��&�h��Y�uw�#6[�ѫ��憃�qxz�p��3���jčj�5] r�?נ�)�K����J!�OM{����Ä	и �~Kj�.��gɜ�Gҋ�|����$<7�q0�%y��$�|�+=~�$�r��֕�*���K���OB��K;!$��ea����)V��p&�q�����f�۔:-݃\����6a�ͷQ+�)Z��:2�LCS7jYA�g0�{���n���J{Gh�Z�ޫ�
�F�Q�;�?�PB7^����obD5D��nBL���5N$ɽ��:�3\�h�\��z�f��=�mAe��GC[H(�y$n�Ō� ikg�ؓC��~N/Mڝ�5#.y1:�'�$gt��<6WE7� |�,O�\]�GM�ҕuaPr3Jm�{�!M����B���F��M[}�X؊�w�\���@-��N������
�Q�3���2TV�����S@h�����-T�L���6�L��D�ua_g�{9�0����.Հ
*�Ak�.B"){7.����1G@�9��Q���2�{%B����Y��y�Q��U\��zP5���^�쀈AW[�4�5��G��	(� �Wu���0I'3���k�_2� �:�N{6Ԯ
�� ee:�}q�����#?��ɝXVv6Z�북��_Q&h�^�ϴ�Jh�	�F2pi[��؊M7�FZ��9�Z:.sV��O�)�ъG��M�]n� L�n�ܝ#/��?�@���!�	2�~����� ����w��P��_Z#C�.�T��4tݏ��cur�nc�7ƿ���d��{��N?�P���5����Z�~�[uqM;$H�T =������9H
��K�qbν�,ToK_��~�,Ȋ�E�>��3�R�U�$	�O���k�(/c�#	¬�Q���)O�!�y��?��Ψb�,�}�h|����=S,b�c-�\���G3�����2U̻�YfU����z�q �χ�6(F]<V��D �g�3:B�����?�1"�����Hl�\�`����/*y[�OɁ4�3���#�^���M��t)����M�Ϯ�p��%7`l���p'�)<�N�MoϺE�Hde��H,.C����fdo�qk�e�7�~���<��m�`��/ eɭ����J�+�M��\��8NF�9������r�JK���+n��N��S"7j��.2�1h��a�����"XV�����������$�|�8W��6�J,\���Y4�+CdE�Y"��5�����]�f_*̥��%��2a�ߑ���@K��5����+�f�Mw]�<k�s`&-5-ڠ��1����D"�B�
�~(nE�(L��[u�J�L@���J�<2΢�?��!�5�A����& ����sU^�+�7�d���u"�.��1\��4B`\3XJ,��)�)u�x<Px���((�͊Z�����`/<����IA� Bm��wEp2� ��T��j�9����]v;�ϐʖd��.�� YӞ[J��il�� �R?F�Nۥ�d9k���p%��jpc�����ZL��on�vT`��@+�x�J({V_E����-�E������|�⛴�P
�**�^נ�_��$sV���9��<���Ɉn�yύ?�*��H勒�m�N)�jX�v�U.MW��ti�g0���Ԫ�,�9x���b�9�˕�o!��;I���g2��=�_ɢ`��l7�F��#�n��,�����O�Tԇ�1��(��8W4֖���Կ��b��� �<"b1#"B�vFd^X8:����_LH
,z�)=.Cq\�V٢u؞�N\wqP�1ՌE����?Qhv��o��J?�'h����%k/����}�%��3� ����;����Q�1R}��q洧U�ͯ�2�e���=c1S	m
�ض�'��<F���U�Y�/U ���ZO�~��'Չn���&���q��
���u�c�x��`���7#*����d���"ңݷX�H�$����|Ze�T��E#��cԺ�9�P�pR����J���n;���]���6X�aþZ'���{�X��e��,�\�c�d�2����oR�O2�?�4`��Ǌ�O�.7��Mx�ꙍ��0�-Ƞ��ɑg(�́���*�ʟ�}���t��ck��>I$���&��L9�(1���(� >A� ����HƧd�l�6���j��}� Y����zJ�v�V��!�����T�����1�͏C�;����\�+����!�o���" �Sf��Q..>-�j/-~����M]R�.WǴ&Y���aA����[m�;\󃱬֛OI!�o
dw,aiR���VU�;�1����,��|-yH!9�$%Niz���+�(������?�N�`����T|)2������#�g1�����73��zB+�.�sd��G��N>TX�>�ߨ�n�{��>eG�,DE��U���m�SN��>���Oy��m�ˑ\p�����ӭ�fq ������_��O�Ʊ�=��Y*5� ��đ��\OU�Sx�h~����֕���ӎ���_<:�<s2y�ͤw�5��S�<�����V�)�%����c�+yY�tK7Vl82�煣����D�H72˙�['��=K�ڙdT*ܰ�DV��eF�J�O���^tf�&EO����m-eo��ґ��~2\��;�i�$�>/��g�k�T�"������/ �ӗm3�����Kp	�W �z���*����w�왿�ά�����	�A����E�Й������@lR;<-�ib��`�w�Wsʹζ���	�LgF3��v�<#��'ߩ�۬_���G�������!����fk޼����C�h��b���H{&@�-�e���#;_3U�[��zՇ�{�)=�����$��5
�]�/��8��������)Ec3��l3O�����W�]�7��I�n����X=�	����	E8�LD��O�����[Y�|Q�ԗJD�$������J[�q&}�A]~��x�ǒQ��#n_»U��u�� �{�h!wԆ���"�\�rߤ4Z��Es�Lu��{l�}^�wu��,���8�W�I'�b\͢�T�~2�Ȍ��9������Q=!�	�f�X��.^<��n���l	�G ed�u���=ǅ�=wO�C������{�o�'�&<3"��C8��?�����v�'z�iϲ�� ��Ŧ�"Ύ�x^�
�T�qBǼ c�-%��}C_��m�t@�8��~P:��`4$s�F��AY/�-k��냪�;�߹� U�����l�Kl���?�9�x��S=��C69|�D�ӊ�wў�0حC��E�:����_ů�����������F�䲭YA�D�^���~���?�j0�6�,4��ܑI�xOe[�`A+�}T?M�o{ڹ�dc�>Ǽ� /�^PF���I�7�7qr���m����VS��}�`m�����1��s��k!O[z���I��3��N~>�ǩO%��@���mg���)�`��"h ~J��Z�$���lj^վ+���b1�7�+�����Yh'�&�^�AEW�k�Rtm��ˁ��+�zn��'?�._ߙ=�*����Ym��/a��e7Mg&D�jk�&��7�G>�6�H!�T,H��t��bѺ#�J��G'[��5�Wn�^u��Y�à�������ZO˅,bs�B+-eI�3������s94v��;�_r�MtM����SBd��#��[�m�5x�{�^����[A�����f����(@�&�v/�ji/>�_ւ��Ӭ`M4�:y_b��_N"�F�:�����D��J��P�_��qn6x	؈�5@6�Q.����; �;�>1�vq�7��[��
c_i �/=c�&�Fx��n?d%���p��R$������x=�����Y�t�iBD)��