��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���,���`�Q �����6�͍	),�6�md|_��n�x�"u������K �5owJh�E��qڑI9����%,%UEwf�x����;.�9��p3��,/�֤����"��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htdʮz_�0�`��@�[D˂8��k�ľF�n�Ԥ��r�τ�u�&&����\l&�$������<H�����}�ƌRS>�(B-~�� ��ڣ�9#M��c��&��C:��pǾE(
'�|�Hۖ4�tgbaY}3�c*����� ����!�_���]̢�X�V����k$bW���5q6耹Q>�װ�����o���/Y�<Ի�C�hQ��N4��K�t�lo�&�2f���2�r�����qgT�Z�Е�~�ΕE(��1ͦǄt�ƕLVE�V�v.��'�=v����h�1A�:,t�3���Quq��N�����=�?�V��a?hgP����d�7[#��l��ۏ/	�:��. �{�˧赂n���ΚI�&�D�u{�"t,�,�`�
V�~���*z`)u�΀/�~��3@�Z#��H#P�!���K����	�?�����:����4�Re�+T��1�ٴp�}�&-kL�D�i/7�M3Η�番	��'M�]����*dE����H�;�f���,�,�B42\���4BE���s@�x�T6`���E?2҂���&��ϡ��K��v�eD��i G�͹Jdo��0�-� \���ӫ���Z [�5��d��዁ԁ5�MM�?p���d�7��½6��%5�Q���	4# Ӗ>�����ĝ��nI����H<��<E�{�D�}����l�3��s	���j~�d��N�0��h�]�7"��~�������\l"�z�ZD����Kd��W�% wTi��8j+l�H�a�"�ypN�����%��J0	s�UVT�w�3��8]V��	�u���p�����/��3��0=	n��
�����aE�cΒ� �xA���[H����+,�2S�����=��1Є0��(�}-^��I�%�n<i�8��f�Z�{{o�}��GhyJ��������4+����5~�l���$-����\��<x�r�($���R��j{!p��A����s�(�)SVz܀�����g�vȾ�Z��f�'ٮ���e�9}:5��/>��[�b�P-��`��[T�;F��c�}� ���������V��Oj�V�+~{Y	�8�!5�����!��(�\�Y.��w�[����� �������r��e���a9h�i�)p�(]�m�� um��_i�5{�?��A�ފ&��{[;�ޯW�1}*B>L��b�.9��ϕ���3A��X�����hӖ���$�Q��՞_�&��cwV�c^r�^X�|����M��#[��y���8�����,�ML�u�E0����=�˂�7�w��*Ia�E��U�Ւ*v���8�M�'�����vz�H�{uݙ�]B>g��@�u�y)��TlTh� ���'�6���E
��p���
ϡwE)�Y���A]�/s������O�2*��W�����Z�["��k����z���yX�|N����",Q ��<Ũ"�"�3����&cZ �Z�m�(�MT�^���G�zG�%��>0������$yXR�u��PC��Rb��u.�Ж���ڴ����3%��Uuh��H��if�א��x:_1�~�(�����v�KUT���h3��`�b��i4�4��_bV��k`�h]��&��.�b�xjbҫ�CP��3�:������[:��Jhk`��� �5|G)e\�wý���w0�@y��ݵ�� �C�H��&x'��:��ˆ���>�ixOd���
#��JzM�.�*��؀���yW'�=WwՖ�Y�J��è3䤙�)!���> jf#�1,S�v�p��-���Aw1���*�O�|�<���RnK�z��A��G��s9:D��f�Ol%�_����T��D�l'{~�S0�F���~۹��_��\HxM���g.���P��X�d�d���*V�3Ht���q���cy�R�	�@��R�����tNv�L{ ���#�U�u{,�Gʍr!�㉥o�Pځ3���h�s�3mK��-+�3#O^+=��u8�򄏼��0ǽ�`?�֋�I�Oۊn
[#_��i�Y��5�Uft���l2��O�BH�Հ��5��,���~4ҎTg���M�Ι���X�4��K���p����[��M�xi=_I|w���I#��w:�����E�÷Z
���
��:>���^���@�osc�Gm�uȗ�Gx�4~��Y|�N��A���zm�\̝ �Q�R�]�m�)-㡀!�9�g��49��ي�JQ����r�����Ȕ�C�<���n�u��6KE���/�>��M��K�5TpD��	�;�%	�7T�\����Q#��5? �2PjqX�iL�E����f��~x�4��$a�������BZlG�	��_������-%=�c��3�)K�����n�]���&=�U����f�]L����eca{@�s��b	�:�\�d�6��"Zd�|��w���$�>[gX �>��<ar�L����ң���MҌ���8���������9�}KT�0�-����m�Z������Y������ua�r�/R YB_���ئ�YwG�U���U�Jt�l���H�V� _��[��{gz�[����v���9_Pz��V��Cゼ�V���$���(Eo�^JI�,�������Πy�<�nl��aB�ޝ��n�Wo�Jn���xI��y����5~x���&-Xp�z�~��d\�8(�!��r5<\�I�>�&Q��_5��S9��+��SJ�َ�5 ���L�1��L�^�T�ޛ�&i�}P"̍�ms� ��yae�@N��Z�bZ�E��wh*�o�!�m��ܻ�ٛ{=Ư������H!���3ȗ�aQ���l�$�	��	ݤ="}������z������0@G��� ZSr��F���>hӼ���Y�:W�v�\��t���P�2��ۑe�&��β_��2#A�W)z�� � Π��w�{���.� kH��"%��va`8��
LEf ��?�{�C^ܪ���l��X���!%�Æ<������b&bW;B��.�zЙ�R�^I,�#O���� u^A����K*�C�+"�)�'w�R����2�Ȧy<\�|�u�^�N�Ӻ,T ��ID���`<���?N%9k����j��8O�0���,�q`_q �S����� '�HY��REr�!��t-]e8pǇ�'Orхc�`��ܴ�5�䗍@��`DS�yu�